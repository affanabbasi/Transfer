magic
tech sky130A
magscale 1 2
timestamp 1607293554
<< nwell >>
rect 10087 7776 21471 7832
rect 29472 7824 42282 7832
rect 50610 7824 63420 7832
rect 29368 7822 42282 7824
rect 50506 7822 63420 7824
rect 28966 7816 42282 7822
rect 50104 7816 63420 7822
rect 26150 7812 42282 7816
rect 47288 7812 63420 7816
rect 23608 7776 42282 7812
rect 44746 7776 63420 7812
rect 10087 4992 63420 7776
rect 10087 4970 21471 4992
rect 23306 4986 42891 4992
rect 23306 4984 24108 4986
rect 26084 4970 42891 4986
rect 44444 4986 63420 4992
rect 44444 4984 45246 4986
rect 47222 4970 63420 4986
rect 16180 4960 18346 4970
rect 26788 4960 28954 4970
rect 37316 4960 39482 4970
rect 47926 4960 50092 4970
rect 58454 4960 60620 4970
<< pwell >>
rect 14268 4282 17364 4286
rect 24876 4282 27972 4286
rect 35404 4282 38500 4286
rect 46014 4282 49110 4286
rect 56542 4282 59638 4286
rect 14268 4272 19740 4282
rect 24876 4272 30348 4282
rect 35404 4272 40876 4282
rect 46014 4272 51486 4282
rect 56542 4272 62014 4282
rect 11870 3860 19740 4272
rect 22478 3860 30348 4272
rect 33006 3860 40876 4272
rect 43616 3860 51486 4272
rect 54144 3860 62014 4272
rect 11870 3850 17364 3860
rect 22478 3850 27972 3860
rect 33006 3850 38500 3860
rect 43616 3850 49110 3860
rect 54144 3850 59638 3860
rect 14268 3846 17364 3850
rect 24876 3846 27972 3850
rect 35404 3846 38500 3850
rect 46014 3846 49110 3850
rect 56542 3846 59638 3850
rect 14279 443 19651 3263
rect 24887 443 30259 3263
rect 35415 443 40787 3263
rect 46025 443 51397 3263
rect 56553 443 61925 3263
<< pmos >>
rect 13560 5205 13960 7205
rect 14018 5205 14418 7205
rect 14476 5205 14876 7205
rect 14934 5205 15334 7205
rect 24168 5205 24568 7205
rect 24626 5205 25026 7205
rect 25084 5205 25484 7205
rect 25542 5205 25942 7205
rect 34696 5205 35096 7205
rect 35154 5205 35554 7205
rect 35612 5205 36012 7205
rect 36070 5205 36470 7205
rect 45306 5205 45706 7205
rect 45764 5205 46164 7205
rect 46222 5205 46622 7205
rect 46680 5205 47080 7205
rect 55834 5205 56234 7205
rect 56292 5205 56692 7205
rect 56750 5205 57150 7205
rect 57208 5205 57608 7205
<< pmoslvt >>
rect 10806 5211 11206 7211
rect 11264 5211 11664 7211
rect 11722 5211 12122 7211
rect 12180 5211 12580 7211
rect 16376 5179 16776 7179
rect 16834 5179 17234 7179
rect 17292 5179 17692 7179
rect 17750 5179 18150 7179
rect 18900 5201 19300 7201
rect 19358 5201 19758 7201
rect 19816 5201 20216 7201
rect 20274 5201 20674 7201
rect 21414 5211 21814 7211
rect 21872 5211 22272 7211
rect 22330 5211 22730 7211
rect 22788 5211 23188 7211
rect 26984 5179 27384 7179
rect 27442 5179 27842 7179
rect 27900 5179 28300 7179
rect 28358 5179 28758 7179
rect 29508 5201 29908 7201
rect 29966 5201 30366 7201
rect 30424 5201 30824 7201
rect 30882 5201 31282 7201
rect 31942 5211 32342 7211
rect 32400 5211 32800 7211
rect 32858 5211 33258 7211
rect 33316 5211 33716 7211
rect 37512 5179 37912 7179
rect 37970 5179 38370 7179
rect 38428 5179 38828 7179
rect 38886 5179 39286 7179
rect 40036 5201 40436 7201
rect 40494 5201 40894 7201
rect 40952 5201 41352 7201
rect 41410 5201 41810 7201
rect 42552 5211 42952 7211
rect 43010 5211 43410 7211
rect 43468 5211 43868 7211
rect 43926 5211 44326 7211
rect 48122 5179 48522 7179
rect 48580 5179 48980 7179
rect 49038 5179 49438 7179
rect 49496 5179 49896 7179
rect 50646 5201 51046 7201
rect 51104 5201 51504 7201
rect 51562 5201 51962 7201
rect 52020 5201 52420 7201
rect 53080 5211 53480 7211
rect 53538 5211 53938 7211
rect 53996 5211 54396 7211
rect 54454 5211 54854 7211
rect 58650 5179 59050 7179
rect 59108 5179 59508 7179
rect 59566 5179 59966 7179
rect 60024 5179 60424 7179
rect 61174 5201 61574 7201
rect 61632 5201 62032 7201
rect 62090 5201 62490 7201
rect 62548 5201 62948 7201
<< nmoslvt >>
rect 12080 4046 14080 4076
rect 17530 4056 19530 4086
rect 22688 4046 24688 4076
rect 28138 4056 30138 4086
rect 33216 4046 35216 4076
rect 38666 4056 40666 4086
rect 43826 4046 45826 4076
rect 49276 4056 51276 4086
rect 54354 4046 56354 4076
rect 59804 4056 61804 4086
rect 14475 653 14875 3053
rect 14933 653 15333 3053
rect 15391 653 15791 3053
rect 15849 653 16249 3053
rect 16307 653 16707 3053
rect 16765 653 17165 3053
rect 17223 653 17623 3053
rect 17681 653 18081 3053
rect 18139 653 18539 3053
rect 18597 653 18997 3053
rect 19055 653 19455 3053
rect 25083 653 25483 3053
rect 25541 653 25941 3053
rect 25999 653 26399 3053
rect 26457 653 26857 3053
rect 26915 653 27315 3053
rect 27373 653 27773 3053
rect 27831 653 28231 3053
rect 28289 653 28689 3053
rect 28747 653 29147 3053
rect 29205 653 29605 3053
rect 29663 653 30063 3053
rect 35611 653 36011 3053
rect 36069 653 36469 3053
rect 36527 653 36927 3053
rect 36985 653 37385 3053
rect 37443 653 37843 3053
rect 37901 653 38301 3053
rect 38359 653 38759 3053
rect 38817 653 39217 3053
rect 39275 653 39675 3053
rect 39733 653 40133 3053
rect 40191 653 40591 3053
rect 46221 653 46621 3053
rect 46679 653 47079 3053
rect 47137 653 47537 3053
rect 47595 653 47995 3053
rect 48053 653 48453 3053
rect 48511 653 48911 3053
rect 48969 653 49369 3053
rect 49427 653 49827 3053
rect 49885 653 50285 3053
rect 50343 653 50743 3053
rect 50801 653 51201 3053
rect 56749 653 57149 3053
rect 57207 653 57607 3053
rect 57665 653 58065 3053
rect 58123 653 58523 3053
rect 58581 653 58981 3053
rect 59039 653 59439 3053
rect 59497 653 59897 3053
rect 59955 653 60355 3053
rect 60413 653 60813 3053
rect 60871 653 61271 3053
rect 61329 653 61729 3053
<< ndiff >>
rect 12080 4122 14080 4134
rect 12080 4088 12092 4122
rect 14068 4088 14080 4122
rect 12080 4076 14080 4088
rect 12080 4034 14080 4046
rect 12080 4000 12092 4034
rect 14068 4000 14080 4034
rect 12080 3988 14080 4000
rect 17530 4132 19530 4144
rect 17530 4098 17542 4132
rect 19518 4098 19530 4132
rect 17530 4086 19530 4098
rect 17530 4044 19530 4056
rect 17530 4010 17542 4044
rect 19518 4010 19530 4044
rect 17530 3998 19530 4010
rect 22688 4122 24688 4134
rect 22688 4088 22700 4122
rect 24676 4088 24688 4122
rect 22688 4076 24688 4088
rect 22688 4034 24688 4046
rect 22688 4000 22700 4034
rect 24676 4000 24688 4034
rect 22688 3988 24688 4000
rect 28138 4132 30138 4144
rect 28138 4098 28150 4132
rect 30126 4098 30138 4132
rect 28138 4086 30138 4098
rect 28138 4044 30138 4056
rect 28138 4010 28150 4044
rect 30126 4010 30138 4044
rect 28138 3998 30138 4010
rect 33216 4122 35216 4134
rect 33216 4088 33228 4122
rect 35204 4088 35216 4122
rect 33216 4076 35216 4088
rect 33216 4034 35216 4046
rect 33216 4000 33228 4034
rect 35204 4000 35216 4034
rect 33216 3988 35216 4000
rect 38666 4132 40666 4144
rect 38666 4098 38678 4132
rect 40654 4098 40666 4132
rect 38666 4086 40666 4098
rect 38666 4044 40666 4056
rect 38666 4010 38678 4044
rect 40654 4010 40666 4044
rect 38666 3998 40666 4010
rect 43826 4122 45826 4134
rect 43826 4088 43838 4122
rect 45814 4088 45826 4122
rect 43826 4076 45826 4088
rect 43826 4034 45826 4046
rect 43826 4000 43838 4034
rect 45814 4000 45826 4034
rect 43826 3988 45826 4000
rect 49276 4132 51276 4144
rect 49276 4098 49288 4132
rect 51264 4098 51276 4132
rect 49276 4086 51276 4098
rect 49276 4044 51276 4056
rect 49276 4010 49288 4044
rect 51264 4010 51276 4044
rect 49276 3998 51276 4010
rect 54354 4122 56354 4134
rect 54354 4088 54366 4122
rect 56342 4088 56354 4122
rect 54354 4076 56354 4088
rect 54354 4034 56354 4046
rect 54354 4000 54366 4034
rect 56342 4000 56354 4034
rect 54354 3988 56354 4000
rect 59804 4132 61804 4144
rect 59804 4098 59816 4132
rect 61792 4098 61804 4132
rect 59804 4086 61804 4098
rect 59804 4044 61804 4056
rect 59804 4010 59816 4044
rect 61792 4010 61804 4044
rect 59804 3998 61804 4010
rect 14417 3041 14475 3053
rect 14417 665 14429 3041
rect 14463 665 14475 3041
rect 14417 653 14475 665
rect 14875 3041 14933 3053
rect 14875 665 14887 3041
rect 14921 665 14933 3041
rect 14875 653 14933 665
rect 15333 3041 15391 3053
rect 15333 665 15345 3041
rect 15379 665 15391 3041
rect 15333 653 15391 665
rect 15791 3041 15849 3053
rect 15791 665 15803 3041
rect 15837 665 15849 3041
rect 15791 653 15849 665
rect 16249 3041 16307 3053
rect 16249 665 16261 3041
rect 16295 665 16307 3041
rect 16249 653 16307 665
rect 16707 3041 16765 3053
rect 16707 665 16719 3041
rect 16753 665 16765 3041
rect 16707 653 16765 665
rect 17165 3041 17223 3053
rect 17165 665 17177 3041
rect 17211 665 17223 3041
rect 17165 653 17223 665
rect 17623 3041 17681 3053
rect 17623 665 17635 3041
rect 17669 665 17681 3041
rect 17623 653 17681 665
rect 18081 3041 18139 3053
rect 18081 665 18093 3041
rect 18127 665 18139 3041
rect 18081 653 18139 665
rect 18539 3041 18597 3053
rect 18539 665 18551 3041
rect 18585 665 18597 3041
rect 18539 653 18597 665
rect 18997 3041 19055 3053
rect 18997 665 19009 3041
rect 19043 665 19055 3041
rect 18997 653 19055 665
rect 19455 3041 19513 3053
rect 19455 665 19467 3041
rect 19501 665 19513 3041
rect 19455 653 19513 665
rect 25025 3041 25083 3053
rect 25025 665 25037 3041
rect 25071 665 25083 3041
rect 25025 653 25083 665
rect 25483 3041 25541 3053
rect 25483 665 25495 3041
rect 25529 665 25541 3041
rect 25483 653 25541 665
rect 25941 3041 25999 3053
rect 25941 665 25953 3041
rect 25987 665 25999 3041
rect 25941 653 25999 665
rect 26399 3041 26457 3053
rect 26399 665 26411 3041
rect 26445 665 26457 3041
rect 26399 653 26457 665
rect 26857 3041 26915 3053
rect 26857 665 26869 3041
rect 26903 665 26915 3041
rect 26857 653 26915 665
rect 27315 3041 27373 3053
rect 27315 665 27327 3041
rect 27361 665 27373 3041
rect 27315 653 27373 665
rect 27773 3041 27831 3053
rect 27773 665 27785 3041
rect 27819 665 27831 3041
rect 27773 653 27831 665
rect 28231 3041 28289 3053
rect 28231 665 28243 3041
rect 28277 665 28289 3041
rect 28231 653 28289 665
rect 28689 3041 28747 3053
rect 28689 665 28701 3041
rect 28735 665 28747 3041
rect 28689 653 28747 665
rect 29147 3041 29205 3053
rect 29147 665 29159 3041
rect 29193 665 29205 3041
rect 29147 653 29205 665
rect 29605 3041 29663 3053
rect 29605 665 29617 3041
rect 29651 665 29663 3041
rect 29605 653 29663 665
rect 30063 3041 30121 3053
rect 30063 665 30075 3041
rect 30109 665 30121 3041
rect 30063 653 30121 665
rect 35553 3041 35611 3053
rect 35553 665 35565 3041
rect 35599 665 35611 3041
rect 35553 653 35611 665
rect 36011 3041 36069 3053
rect 36011 665 36023 3041
rect 36057 665 36069 3041
rect 36011 653 36069 665
rect 36469 3041 36527 3053
rect 36469 665 36481 3041
rect 36515 665 36527 3041
rect 36469 653 36527 665
rect 36927 3041 36985 3053
rect 36927 665 36939 3041
rect 36973 665 36985 3041
rect 36927 653 36985 665
rect 37385 3041 37443 3053
rect 37385 665 37397 3041
rect 37431 665 37443 3041
rect 37385 653 37443 665
rect 37843 3041 37901 3053
rect 37843 665 37855 3041
rect 37889 665 37901 3041
rect 37843 653 37901 665
rect 38301 3041 38359 3053
rect 38301 665 38313 3041
rect 38347 665 38359 3041
rect 38301 653 38359 665
rect 38759 3041 38817 3053
rect 38759 665 38771 3041
rect 38805 665 38817 3041
rect 38759 653 38817 665
rect 39217 3041 39275 3053
rect 39217 665 39229 3041
rect 39263 665 39275 3041
rect 39217 653 39275 665
rect 39675 3041 39733 3053
rect 39675 665 39687 3041
rect 39721 665 39733 3041
rect 39675 653 39733 665
rect 40133 3041 40191 3053
rect 40133 665 40145 3041
rect 40179 665 40191 3041
rect 40133 653 40191 665
rect 40591 3041 40649 3053
rect 40591 665 40603 3041
rect 40637 665 40649 3041
rect 40591 653 40649 665
rect 46163 3041 46221 3053
rect 46163 665 46175 3041
rect 46209 665 46221 3041
rect 46163 653 46221 665
rect 46621 3041 46679 3053
rect 46621 665 46633 3041
rect 46667 665 46679 3041
rect 46621 653 46679 665
rect 47079 3041 47137 3053
rect 47079 665 47091 3041
rect 47125 665 47137 3041
rect 47079 653 47137 665
rect 47537 3041 47595 3053
rect 47537 665 47549 3041
rect 47583 665 47595 3041
rect 47537 653 47595 665
rect 47995 3041 48053 3053
rect 47995 665 48007 3041
rect 48041 665 48053 3041
rect 47995 653 48053 665
rect 48453 3041 48511 3053
rect 48453 665 48465 3041
rect 48499 665 48511 3041
rect 48453 653 48511 665
rect 48911 3041 48969 3053
rect 48911 665 48923 3041
rect 48957 665 48969 3041
rect 48911 653 48969 665
rect 49369 3041 49427 3053
rect 49369 665 49381 3041
rect 49415 665 49427 3041
rect 49369 653 49427 665
rect 49827 3041 49885 3053
rect 49827 665 49839 3041
rect 49873 665 49885 3041
rect 49827 653 49885 665
rect 50285 3041 50343 3053
rect 50285 665 50297 3041
rect 50331 665 50343 3041
rect 50285 653 50343 665
rect 50743 3041 50801 3053
rect 50743 665 50755 3041
rect 50789 665 50801 3041
rect 50743 653 50801 665
rect 51201 3041 51259 3053
rect 51201 665 51213 3041
rect 51247 665 51259 3041
rect 51201 653 51259 665
rect 56691 3041 56749 3053
rect 56691 665 56703 3041
rect 56737 665 56749 3041
rect 56691 653 56749 665
rect 57149 3041 57207 3053
rect 57149 665 57161 3041
rect 57195 665 57207 3041
rect 57149 653 57207 665
rect 57607 3041 57665 3053
rect 57607 665 57619 3041
rect 57653 665 57665 3041
rect 57607 653 57665 665
rect 58065 3041 58123 3053
rect 58065 665 58077 3041
rect 58111 665 58123 3041
rect 58065 653 58123 665
rect 58523 3041 58581 3053
rect 58523 665 58535 3041
rect 58569 665 58581 3041
rect 58523 653 58581 665
rect 58981 3041 59039 3053
rect 58981 665 58993 3041
rect 59027 665 59039 3041
rect 58981 653 59039 665
rect 59439 3041 59497 3053
rect 59439 665 59451 3041
rect 59485 665 59497 3041
rect 59439 653 59497 665
rect 59897 3041 59955 3053
rect 59897 665 59909 3041
rect 59943 665 59955 3041
rect 59897 653 59955 665
rect 60355 3041 60413 3053
rect 60355 665 60367 3041
rect 60401 665 60413 3041
rect 60355 653 60413 665
rect 60813 3041 60871 3053
rect 60813 665 60825 3041
rect 60859 665 60871 3041
rect 60813 653 60871 665
rect 61271 3041 61329 3053
rect 61271 665 61283 3041
rect 61317 665 61329 3041
rect 61271 653 61329 665
rect 61729 3041 61787 3053
rect 61729 665 61741 3041
rect 61775 665 61787 3041
rect 61729 653 61787 665
<< pdiff >>
rect 10748 7199 10806 7211
rect 10748 5223 10760 7199
rect 10794 5223 10806 7199
rect 10748 5211 10806 5223
rect 11206 7199 11264 7211
rect 11206 5223 11218 7199
rect 11252 5223 11264 7199
rect 11206 5211 11264 5223
rect 11664 7199 11722 7211
rect 11664 5223 11676 7199
rect 11710 5223 11722 7199
rect 11664 5211 11722 5223
rect 12122 7199 12180 7211
rect 12122 5223 12134 7199
rect 12168 5223 12180 7199
rect 12122 5211 12180 5223
rect 12580 7199 12638 7211
rect 12580 5223 12592 7199
rect 12626 5223 12638 7199
rect 12580 5211 12638 5223
rect 13502 7193 13560 7205
rect 13502 5217 13514 7193
rect 13548 5217 13560 7193
rect 13502 5205 13560 5217
rect 13960 7193 14018 7205
rect 13960 5217 13972 7193
rect 14006 5217 14018 7193
rect 13960 5205 14018 5217
rect 14418 7193 14476 7205
rect 14418 5217 14430 7193
rect 14464 5217 14476 7193
rect 14418 5205 14476 5217
rect 14876 7193 14934 7205
rect 14876 5217 14888 7193
rect 14922 5217 14934 7193
rect 14876 5205 14934 5217
rect 15334 7193 15392 7205
rect 15334 5217 15346 7193
rect 15380 5217 15392 7193
rect 15334 5205 15392 5217
rect 16318 7167 16376 7179
rect 16318 5191 16330 7167
rect 16364 5191 16376 7167
rect 16318 5179 16376 5191
rect 16776 7167 16834 7179
rect 16776 5191 16788 7167
rect 16822 5191 16834 7167
rect 16776 5179 16834 5191
rect 17234 7167 17292 7179
rect 17234 5191 17246 7167
rect 17280 5191 17292 7167
rect 17234 5179 17292 5191
rect 17692 7167 17750 7179
rect 17692 5191 17704 7167
rect 17738 5191 17750 7167
rect 17692 5179 17750 5191
rect 18150 7167 18208 7179
rect 18150 5191 18162 7167
rect 18196 5191 18208 7167
rect 18150 5179 18208 5191
rect 18842 7189 18900 7201
rect 18842 5213 18854 7189
rect 18888 5213 18900 7189
rect 18842 5201 18900 5213
rect 19300 7189 19358 7201
rect 19300 5213 19312 7189
rect 19346 5213 19358 7189
rect 19300 5201 19358 5213
rect 19758 7189 19816 7201
rect 19758 5213 19770 7189
rect 19804 5213 19816 7189
rect 19758 5201 19816 5213
rect 20216 7189 20274 7201
rect 20216 5213 20228 7189
rect 20262 5213 20274 7189
rect 20216 5201 20274 5213
rect 20674 7189 20732 7201
rect 20674 5213 20686 7189
rect 20720 5213 20732 7189
rect 20674 5201 20732 5213
rect 21356 7199 21414 7211
rect 21356 5223 21368 7199
rect 21402 5223 21414 7199
rect 21356 5211 21414 5223
rect 21814 7199 21872 7211
rect 21814 5223 21826 7199
rect 21860 5223 21872 7199
rect 21814 5211 21872 5223
rect 22272 7199 22330 7211
rect 22272 5223 22284 7199
rect 22318 5223 22330 7199
rect 22272 5211 22330 5223
rect 22730 7199 22788 7211
rect 22730 5223 22742 7199
rect 22776 5223 22788 7199
rect 22730 5211 22788 5223
rect 23188 7199 23246 7211
rect 23188 5223 23200 7199
rect 23234 5223 23246 7199
rect 23188 5211 23246 5223
rect 24110 7193 24168 7205
rect 24110 5217 24122 7193
rect 24156 5217 24168 7193
rect 24110 5205 24168 5217
rect 24568 7193 24626 7205
rect 24568 5217 24580 7193
rect 24614 5217 24626 7193
rect 24568 5205 24626 5217
rect 25026 7193 25084 7205
rect 25026 5217 25038 7193
rect 25072 5217 25084 7193
rect 25026 5205 25084 5217
rect 25484 7193 25542 7205
rect 25484 5217 25496 7193
rect 25530 5217 25542 7193
rect 25484 5205 25542 5217
rect 25942 7193 26000 7205
rect 25942 5217 25954 7193
rect 25988 5217 26000 7193
rect 25942 5205 26000 5217
rect 26926 7167 26984 7179
rect 26926 5191 26938 7167
rect 26972 5191 26984 7167
rect 26926 5179 26984 5191
rect 27384 7167 27442 7179
rect 27384 5191 27396 7167
rect 27430 5191 27442 7167
rect 27384 5179 27442 5191
rect 27842 7167 27900 7179
rect 27842 5191 27854 7167
rect 27888 5191 27900 7167
rect 27842 5179 27900 5191
rect 28300 7167 28358 7179
rect 28300 5191 28312 7167
rect 28346 5191 28358 7167
rect 28300 5179 28358 5191
rect 28758 7167 28816 7179
rect 28758 5191 28770 7167
rect 28804 5191 28816 7167
rect 28758 5179 28816 5191
rect 29450 7189 29508 7201
rect 29450 5213 29462 7189
rect 29496 5213 29508 7189
rect 29450 5201 29508 5213
rect 29908 7189 29966 7201
rect 29908 5213 29920 7189
rect 29954 5213 29966 7189
rect 29908 5201 29966 5213
rect 30366 7189 30424 7201
rect 30366 5213 30378 7189
rect 30412 5213 30424 7189
rect 30366 5201 30424 5213
rect 30824 7189 30882 7201
rect 30824 5213 30836 7189
rect 30870 5213 30882 7189
rect 30824 5201 30882 5213
rect 31282 7189 31340 7201
rect 31282 5213 31294 7189
rect 31328 5213 31340 7189
rect 31282 5201 31340 5213
rect 31884 7199 31942 7211
rect 31884 5223 31896 7199
rect 31930 5223 31942 7199
rect 31884 5211 31942 5223
rect 32342 7199 32400 7211
rect 32342 5223 32354 7199
rect 32388 5223 32400 7199
rect 32342 5211 32400 5223
rect 32800 7199 32858 7211
rect 32800 5223 32812 7199
rect 32846 5223 32858 7199
rect 32800 5211 32858 5223
rect 33258 7199 33316 7211
rect 33258 5223 33270 7199
rect 33304 5223 33316 7199
rect 33258 5211 33316 5223
rect 33716 7199 33774 7211
rect 33716 5223 33728 7199
rect 33762 5223 33774 7199
rect 33716 5211 33774 5223
rect 34638 7193 34696 7205
rect 34638 5217 34650 7193
rect 34684 5217 34696 7193
rect 34638 5205 34696 5217
rect 35096 7193 35154 7205
rect 35096 5217 35108 7193
rect 35142 5217 35154 7193
rect 35096 5205 35154 5217
rect 35554 7193 35612 7205
rect 35554 5217 35566 7193
rect 35600 5217 35612 7193
rect 35554 5205 35612 5217
rect 36012 7193 36070 7205
rect 36012 5217 36024 7193
rect 36058 5217 36070 7193
rect 36012 5205 36070 5217
rect 36470 7193 36528 7205
rect 36470 5217 36482 7193
rect 36516 5217 36528 7193
rect 36470 5205 36528 5217
rect 37454 7167 37512 7179
rect 37454 5191 37466 7167
rect 37500 5191 37512 7167
rect 37454 5179 37512 5191
rect 37912 7167 37970 7179
rect 37912 5191 37924 7167
rect 37958 5191 37970 7167
rect 37912 5179 37970 5191
rect 38370 7167 38428 7179
rect 38370 5191 38382 7167
rect 38416 5191 38428 7167
rect 38370 5179 38428 5191
rect 38828 7167 38886 7179
rect 38828 5191 38840 7167
rect 38874 5191 38886 7167
rect 38828 5179 38886 5191
rect 39286 7167 39344 7179
rect 39286 5191 39298 7167
rect 39332 5191 39344 7167
rect 39286 5179 39344 5191
rect 39978 7189 40036 7201
rect 39978 5213 39990 7189
rect 40024 5213 40036 7189
rect 39978 5201 40036 5213
rect 40436 7189 40494 7201
rect 40436 5213 40448 7189
rect 40482 5213 40494 7189
rect 40436 5201 40494 5213
rect 40894 7189 40952 7201
rect 40894 5213 40906 7189
rect 40940 5213 40952 7189
rect 40894 5201 40952 5213
rect 41352 7189 41410 7201
rect 41352 5213 41364 7189
rect 41398 5213 41410 7189
rect 41352 5201 41410 5213
rect 41810 7189 41868 7201
rect 41810 5213 41822 7189
rect 41856 5213 41868 7189
rect 41810 5201 41868 5213
rect 42494 7199 42552 7211
rect 42494 5223 42506 7199
rect 42540 5223 42552 7199
rect 42494 5211 42552 5223
rect 42952 7199 43010 7211
rect 42952 5223 42964 7199
rect 42998 5223 43010 7199
rect 42952 5211 43010 5223
rect 43410 7199 43468 7211
rect 43410 5223 43422 7199
rect 43456 5223 43468 7199
rect 43410 5211 43468 5223
rect 43868 7199 43926 7211
rect 43868 5223 43880 7199
rect 43914 5223 43926 7199
rect 43868 5211 43926 5223
rect 44326 7199 44384 7211
rect 44326 5223 44338 7199
rect 44372 5223 44384 7199
rect 44326 5211 44384 5223
rect 45248 7193 45306 7205
rect 45248 5217 45260 7193
rect 45294 5217 45306 7193
rect 45248 5205 45306 5217
rect 45706 7193 45764 7205
rect 45706 5217 45718 7193
rect 45752 5217 45764 7193
rect 45706 5205 45764 5217
rect 46164 7193 46222 7205
rect 46164 5217 46176 7193
rect 46210 5217 46222 7193
rect 46164 5205 46222 5217
rect 46622 7193 46680 7205
rect 46622 5217 46634 7193
rect 46668 5217 46680 7193
rect 46622 5205 46680 5217
rect 47080 7193 47138 7205
rect 47080 5217 47092 7193
rect 47126 5217 47138 7193
rect 47080 5205 47138 5217
rect 48064 7167 48122 7179
rect 48064 5191 48076 7167
rect 48110 5191 48122 7167
rect 48064 5179 48122 5191
rect 48522 7167 48580 7179
rect 48522 5191 48534 7167
rect 48568 5191 48580 7167
rect 48522 5179 48580 5191
rect 48980 7167 49038 7179
rect 48980 5191 48992 7167
rect 49026 5191 49038 7167
rect 48980 5179 49038 5191
rect 49438 7167 49496 7179
rect 49438 5191 49450 7167
rect 49484 5191 49496 7167
rect 49438 5179 49496 5191
rect 49896 7167 49954 7179
rect 49896 5191 49908 7167
rect 49942 5191 49954 7167
rect 49896 5179 49954 5191
rect 50588 7189 50646 7201
rect 50588 5213 50600 7189
rect 50634 5213 50646 7189
rect 50588 5201 50646 5213
rect 51046 7189 51104 7201
rect 51046 5213 51058 7189
rect 51092 5213 51104 7189
rect 51046 5201 51104 5213
rect 51504 7189 51562 7201
rect 51504 5213 51516 7189
rect 51550 5213 51562 7189
rect 51504 5201 51562 5213
rect 51962 7189 52020 7201
rect 51962 5213 51974 7189
rect 52008 5213 52020 7189
rect 51962 5201 52020 5213
rect 52420 7189 52478 7201
rect 52420 5213 52432 7189
rect 52466 5213 52478 7189
rect 52420 5201 52478 5213
rect 53022 7199 53080 7211
rect 53022 5223 53034 7199
rect 53068 5223 53080 7199
rect 53022 5211 53080 5223
rect 53480 7199 53538 7211
rect 53480 5223 53492 7199
rect 53526 5223 53538 7199
rect 53480 5211 53538 5223
rect 53938 7199 53996 7211
rect 53938 5223 53950 7199
rect 53984 5223 53996 7199
rect 53938 5211 53996 5223
rect 54396 7199 54454 7211
rect 54396 5223 54408 7199
rect 54442 5223 54454 7199
rect 54396 5211 54454 5223
rect 54854 7199 54912 7211
rect 54854 5223 54866 7199
rect 54900 5223 54912 7199
rect 54854 5211 54912 5223
rect 55776 7193 55834 7205
rect 55776 5217 55788 7193
rect 55822 5217 55834 7193
rect 55776 5205 55834 5217
rect 56234 7193 56292 7205
rect 56234 5217 56246 7193
rect 56280 5217 56292 7193
rect 56234 5205 56292 5217
rect 56692 7193 56750 7205
rect 56692 5217 56704 7193
rect 56738 5217 56750 7193
rect 56692 5205 56750 5217
rect 57150 7193 57208 7205
rect 57150 5217 57162 7193
rect 57196 5217 57208 7193
rect 57150 5205 57208 5217
rect 57608 7193 57666 7205
rect 57608 5217 57620 7193
rect 57654 5217 57666 7193
rect 57608 5205 57666 5217
rect 58592 7167 58650 7179
rect 58592 5191 58604 7167
rect 58638 5191 58650 7167
rect 58592 5179 58650 5191
rect 59050 7167 59108 7179
rect 59050 5191 59062 7167
rect 59096 5191 59108 7167
rect 59050 5179 59108 5191
rect 59508 7167 59566 7179
rect 59508 5191 59520 7167
rect 59554 5191 59566 7167
rect 59508 5179 59566 5191
rect 59966 7167 60024 7179
rect 59966 5191 59978 7167
rect 60012 5191 60024 7167
rect 59966 5179 60024 5191
rect 60424 7167 60482 7179
rect 60424 5191 60436 7167
rect 60470 5191 60482 7167
rect 60424 5179 60482 5191
rect 61116 7189 61174 7201
rect 61116 5213 61128 7189
rect 61162 5213 61174 7189
rect 61116 5201 61174 5213
rect 61574 7189 61632 7201
rect 61574 5213 61586 7189
rect 61620 5213 61632 7189
rect 61574 5201 61632 5213
rect 62032 7189 62090 7201
rect 62032 5213 62044 7189
rect 62078 5213 62090 7189
rect 62032 5201 62090 5213
rect 62490 7189 62548 7201
rect 62490 5213 62502 7189
rect 62536 5213 62548 7189
rect 62490 5201 62548 5213
rect 62948 7189 63006 7201
rect 62948 5213 62960 7189
rect 62994 5213 63006 7189
rect 62948 5201 63006 5213
<< ndiffc >>
rect 12092 4088 14068 4122
rect 12092 4000 14068 4034
rect 17542 4098 19518 4132
rect 17542 4010 19518 4044
rect 22700 4088 24676 4122
rect 22700 4000 24676 4034
rect 28150 4098 30126 4132
rect 28150 4010 30126 4044
rect 33228 4088 35204 4122
rect 33228 4000 35204 4034
rect 38678 4098 40654 4132
rect 38678 4010 40654 4044
rect 43838 4088 45814 4122
rect 43838 4000 45814 4034
rect 49288 4098 51264 4132
rect 49288 4010 51264 4044
rect 54366 4088 56342 4122
rect 54366 4000 56342 4034
rect 59816 4098 61792 4132
rect 59816 4010 61792 4044
rect 14429 665 14463 3041
rect 14887 665 14921 3041
rect 15345 665 15379 3041
rect 15803 665 15837 3041
rect 16261 665 16295 3041
rect 16719 665 16753 3041
rect 17177 665 17211 3041
rect 17635 665 17669 3041
rect 18093 665 18127 3041
rect 18551 665 18585 3041
rect 19009 665 19043 3041
rect 19467 665 19501 3041
rect 25037 665 25071 3041
rect 25495 665 25529 3041
rect 25953 665 25987 3041
rect 26411 665 26445 3041
rect 26869 665 26903 3041
rect 27327 665 27361 3041
rect 27785 665 27819 3041
rect 28243 665 28277 3041
rect 28701 665 28735 3041
rect 29159 665 29193 3041
rect 29617 665 29651 3041
rect 30075 665 30109 3041
rect 35565 665 35599 3041
rect 36023 665 36057 3041
rect 36481 665 36515 3041
rect 36939 665 36973 3041
rect 37397 665 37431 3041
rect 37855 665 37889 3041
rect 38313 665 38347 3041
rect 38771 665 38805 3041
rect 39229 665 39263 3041
rect 39687 665 39721 3041
rect 40145 665 40179 3041
rect 40603 665 40637 3041
rect 46175 665 46209 3041
rect 46633 665 46667 3041
rect 47091 665 47125 3041
rect 47549 665 47583 3041
rect 48007 665 48041 3041
rect 48465 665 48499 3041
rect 48923 665 48957 3041
rect 49381 665 49415 3041
rect 49839 665 49873 3041
rect 50297 665 50331 3041
rect 50755 665 50789 3041
rect 51213 665 51247 3041
rect 56703 665 56737 3041
rect 57161 665 57195 3041
rect 57619 665 57653 3041
rect 58077 665 58111 3041
rect 58535 665 58569 3041
rect 58993 665 59027 3041
rect 59451 665 59485 3041
rect 59909 665 59943 3041
rect 60367 665 60401 3041
rect 60825 665 60859 3041
rect 61283 665 61317 3041
rect 61741 665 61775 3041
<< pdiffc >>
rect 10760 5223 10794 7199
rect 11218 5223 11252 7199
rect 11676 5223 11710 7199
rect 12134 5223 12168 7199
rect 12592 5223 12626 7199
rect 13514 5217 13548 7193
rect 13972 5217 14006 7193
rect 14430 5217 14464 7193
rect 14888 5217 14922 7193
rect 15346 5217 15380 7193
rect 16330 5191 16364 7167
rect 16788 5191 16822 7167
rect 17246 5191 17280 7167
rect 17704 5191 17738 7167
rect 18162 5191 18196 7167
rect 18854 5213 18888 7189
rect 19312 5213 19346 7189
rect 19770 5213 19804 7189
rect 20228 5213 20262 7189
rect 20686 5213 20720 7189
rect 21368 5223 21402 7199
rect 21826 5223 21860 7199
rect 22284 5223 22318 7199
rect 22742 5223 22776 7199
rect 23200 5223 23234 7199
rect 24122 5217 24156 7193
rect 24580 5217 24614 7193
rect 25038 5217 25072 7193
rect 25496 5217 25530 7193
rect 25954 5217 25988 7193
rect 26938 5191 26972 7167
rect 27396 5191 27430 7167
rect 27854 5191 27888 7167
rect 28312 5191 28346 7167
rect 28770 5191 28804 7167
rect 29462 5213 29496 7189
rect 29920 5213 29954 7189
rect 30378 5213 30412 7189
rect 30836 5213 30870 7189
rect 31294 5213 31328 7189
rect 31896 5223 31930 7199
rect 32354 5223 32388 7199
rect 32812 5223 32846 7199
rect 33270 5223 33304 7199
rect 33728 5223 33762 7199
rect 34650 5217 34684 7193
rect 35108 5217 35142 7193
rect 35566 5217 35600 7193
rect 36024 5217 36058 7193
rect 36482 5217 36516 7193
rect 37466 5191 37500 7167
rect 37924 5191 37958 7167
rect 38382 5191 38416 7167
rect 38840 5191 38874 7167
rect 39298 5191 39332 7167
rect 39990 5213 40024 7189
rect 40448 5213 40482 7189
rect 40906 5213 40940 7189
rect 41364 5213 41398 7189
rect 41822 5213 41856 7189
rect 42506 5223 42540 7199
rect 42964 5223 42998 7199
rect 43422 5223 43456 7199
rect 43880 5223 43914 7199
rect 44338 5223 44372 7199
rect 45260 5217 45294 7193
rect 45718 5217 45752 7193
rect 46176 5217 46210 7193
rect 46634 5217 46668 7193
rect 47092 5217 47126 7193
rect 48076 5191 48110 7167
rect 48534 5191 48568 7167
rect 48992 5191 49026 7167
rect 49450 5191 49484 7167
rect 49908 5191 49942 7167
rect 50600 5213 50634 7189
rect 51058 5213 51092 7189
rect 51516 5213 51550 7189
rect 51974 5213 52008 7189
rect 52432 5213 52466 7189
rect 53034 5223 53068 7199
rect 53492 5223 53526 7199
rect 53950 5223 53984 7199
rect 54408 5223 54442 7199
rect 54866 5223 54900 7199
rect 55788 5217 55822 7193
rect 56246 5217 56280 7193
rect 56704 5217 56738 7193
rect 57162 5217 57196 7193
rect 57620 5217 57654 7193
rect 58604 5191 58638 7167
rect 59062 5191 59096 7167
rect 59520 5191 59554 7167
rect 59978 5191 60012 7167
rect 60436 5191 60470 7167
rect 61128 5213 61162 7189
rect 61586 5213 61620 7189
rect 62044 5213 62078 7189
rect 62502 5213 62536 7189
rect 62960 5213 62994 7189
<< psubdiff >>
rect 11906 4202 12002 4236
rect 14158 4202 14254 4236
rect 11906 4140 11940 4202
rect 14220 4140 14254 4202
rect 11906 3920 11940 3982
rect 14220 3920 14254 3982
rect 11906 3886 12002 3920
rect 14158 3886 14254 3920
rect 17356 4212 17452 4246
rect 19608 4212 19704 4246
rect 17356 4150 17390 4212
rect 19670 4150 19704 4212
rect 17356 3930 17390 3992
rect 19670 3930 19704 3992
rect 17356 3896 17452 3930
rect 19608 3896 19704 3930
rect 22514 4202 22610 4236
rect 24766 4202 24862 4236
rect 22514 4140 22548 4202
rect 24828 4140 24862 4202
rect 22514 3920 22548 3982
rect 24828 3920 24862 3982
rect 22514 3886 22610 3920
rect 24766 3886 24862 3920
rect 27964 4212 28060 4246
rect 30216 4212 30312 4246
rect 27964 4150 27998 4212
rect 30278 4150 30312 4212
rect 27964 3930 27998 3992
rect 30278 3930 30312 3992
rect 27964 3896 28060 3930
rect 30216 3896 30312 3930
rect 33042 4202 33138 4236
rect 35294 4202 35390 4236
rect 33042 4140 33076 4202
rect 35356 4140 35390 4202
rect 33042 3920 33076 3982
rect 35356 3920 35390 3982
rect 33042 3886 33138 3920
rect 35294 3886 35390 3920
rect 38492 4212 38588 4246
rect 40744 4212 40840 4246
rect 38492 4150 38526 4212
rect 40806 4150 40840 4212
rect 38492 3930 38526 3992
rect 40806 3930 40840 3992
rect 38492 3896 38588 3930
rect 40744 3896 40840 3930
rect 43652 4202 43748 4236
rect 45904 4202 46000 4236
rect 43652 4140 43686 4202
rect 45966 4140 46000 4202
rect 43652 3920 43686 3982
rect 45966 3920 46000 3982
rect 43652 3886 43748 3920
rect 45904 3886 46000 3920
rect 49102 4212 49198 4246
rect 51354 4212 51450 4246
rect 49102 4150 49136 4212
rect 51416 4150 51450 4212
rect 49102 3930 49136 3992
rect 51416 3930 51450 3992
rect 49102 3896 49198 3930
rect 51354 3896 51450 3930
rect 54180 4202 54276 4236
rect 56432 4202 56528 4236
rect 54180 4140 54214 4202
rect 56494 4140 56528 4202
rect 54180 3920 54214 3982
rect 56494 3920 56528 3982
rect 54180 3886 54276 3920
rect 56432 3886 56528 3920
rect 59630 4212 59726 4246
rect 61882 4212 61978 4246
rect 59630 4150 59664 4212
rect 61944 4150 61978 4212
rect 59630 3930 59664 3992
rect 61944 3930 61978 3992
rect 59630 3896 59726 3930
rect 61882 3896 61978 3930
rect 14315 3193 14411 3227
rect 19519 3193 19615 3227
rect 14315 3131 14349 3193
rect 19581 3131 19615 3193
rect 14315 513 14349 575
rect 19581 513 19615 575
rect 14315 479 14411 513
rect 19519 479 19615 513
rect 24923 3193 25019 3227
rect 30127 3193 30223 3227
rect 24923 3131 24957 3193
rect 30189 3131 30223 3193
rect 24923 513 24957 575
rect 30189 513 30223 575
rect 24923 479 25019 513
rect 30127 479 30223 513
rect 35451 3193 35547 3227
rect 40655 3193 40751 3227
rect 35451 3131 35485 3193
rect 40717 3131 40751 3193
rect 35451 513 35485 575
rect 40717 513 40751 575
rect 35451 479 35547 513
rect 40655 479 40751 513
rect 46061 3193 46157 3227
rect 51265 3193 51361 3227
rect 46061 3131 46095 3193
rect 51327 3131 51361 3193
rect 46061 513 46095 575
rect 51327 513 51361 575
rect 46061 479 46157 513
rect 51265 479 51361 513
rect 56589 3193 56685 3227
rect 61793 3193 61889 3227
rect 56589 3131 56623 3193
rect 61855 3131 61889 3193
rect 56589 513 56623 575
rect 61855 513 61889 575
rect 56589 479 56685 513
rect 61793 479 61889 513
rect 14244 268 19776 322
rect 14244 264 18590 268
rect 14244 258 15722 264
rect 14244 142 14828 258
rect 14986 148 15722 258
rect 15880 148 17492 264
rect 17650 152 18590 264
rect 18748 152 19776 268
rect 17650 148 19776 152
rect 14986 142 19776 148
rect 14244 94 19776 142
rect 24852 268 30384 322
rect 24852 264 29198 268
rect 24852 258 26330 264
rect 24852 142 25436 258
rect 25594 148 26330 258
rect 26488 148 28100 264
rect 28258 152 29198 264
rect 29356 152 30384 268
rect 28258 148 30384 152
rect 25594 142 30384 148
rect 24852 94 30384 142
rect 35380 268 40912 322
rect 35380 264 39726 268
rect 35380 258 36858 264
rect 35380 142 35964 258
rect 36122 148 36858 258
rect 37016 148 38628 264
rect 38786 152 39726 264
rect 39884 152 40912 268
rect 38786 148 40912 152
rect 36122 142 40912 148
rect 35380 94 40912 142
rect 45990 268 51522 322
rect 45990 264 50336 268
rect 45990 258 47468 264
rect 45990 142 46574 258
rect 46732 148 47468 258
rect 47626 148 49238 264
rect 49396 152 50336 264
rect 50494 152 51522 268
rect 49396 148 51522 152
rect 46732 142 51522 148
rect 45990 94 51522 142
rect 56518 268 62050 322
rect 56518 264 60864 268
rect 56518 258 57996 264
rect 56518 142 57102 258
rect 57260 148 57996 258
rect 58154 148 59766 264
rect 59924 152 60864 264
rect 61022 152 62050 268
rect 59924 148 62050 152
rect 57260 142 62050 148
rect 56518 94 62050 142
<< nsubdiff >>
rect 18416 7710 20886 7730
rect 29024 7710 31494 7730
rect 39552 7710 42022 7730
rect 50162 7710 52632 7730
rect 60690 7710 63160 7730
rect 15422 7708 20886 7710
rect 26030 7708 31494 7710
rect 36558 7708 42022 7710
rect 47168 7708 52632 7710
rect 57696 7708 63160 7710
rect 10658 7696 20886 7708
rect 10658 7678 16708 7696
rect 10658 7668 13916 7678
rect 10658 7658 12074 7668
rect 10658 7564 11140 7658
rect 11276 7574 12074 7658
rect 12210 7588 13916 7668
rect 14028 7670 16708 7678
rect 14028 7588 14834 7670
rect 12210 7580 14834 7588
rect 14946 7594 16708 7670
rect 16814 7690 20886 7696
rect 16814 7594 17670 7690
rect 14946 7588 17670 7594
rect 17776 7684 20886 7690
rect 17776 7682 20194 7684
rect 17776 7590 19248 7682
rect 19338 7592 20194 7682
rect 20284 7592 20886 7684
rect 19338 7590 20886 7592
rect 17776 7588 20886 7590
rect 14946 7580 20886 7588
rect 12210 7574 20886 7580
rect 11276 7564 20886 7574
rect 10658 7556 20886 7564
rect 10658 7548 12780 7556
rect 15422 7552 20886 7556
rect 18416 7548 20886 7552
rect 21266 7696 31494 7708
rect 21266 7678 27316 7696
rect 21266 7668 24524 7678
rect 21266 7658 22682 7668
rect 21266 7564 21748 7658
rect 21884 7574 22682 7658
rect 22818 7588 24524 7668
rect 24636 7670 27316 7678
rect 24636 7588 25442 7670
rect 22818 7580 25442 7588
rect 25554 7594 27316 7670
rect 27422 7690 31494 7696
rect 27422 7594 28278 7690
rect 25554 7588 28278 7594
rect 28384 7684 31494 7690
rect 28384 7682 30802 7684
rect 28384 7590 29856 7682
rect 29946 7592 30802 7682
rect 30892 7592 31494 7684
rect 29946 7590 31494 7592
rect 28384 7588 31494 7590
rect 25554 7580 31494 7588
rect 22818 7574 31494 7580
rect 21884 7564 31494 7574
rect 21266 7556 31494 7564
rect 21266 7548 23388 7556
rect 26030 7552 31494 7556
rect 29024 7548 31494 7552
rect 31794 7696 42022 7708
rect 31794 7678 37844 7696
rect 31794 7668 35052 7678
rect 31794 7658 33210 7668
rect 31794 7564 32276 7658
rect 32412 7574 33210 7658
rect 33346 7588 35052 7668
rect 35164 7670 37844 7678
rect 35164 7588 35970 7670
rect 33346 7580 35970 7588
rect 36082 7594 37844 7670
rect 37950 7690 42022 7696
rect 37950 7594 38806 7690
rect 36082 7588 38806 7594
rect 38912 7684 42022 7690
rect 38912 7682 41330 7684
rect 38912 7590 40384 7682
rect 40474 7592 41330 7682
rect 41420 7592 42022 7684
rect 40474 7590 42022 7592
rect 38912 7588 42022 7590
rect 36082 7580 42022 7588
rect 33346 7574 42022 7580
rect 32412 7564 42022 7574
rect 31794 7556 42022 7564
rect 31794 7548 33916 7556
rect 36558 7552 42022 7556
rect 39552 7548 42022 7552
rect 42404 7696 52632 7708
rect 42404 7678 48454 7696
rect 42404 7668 45662 7678
rect 42404 7658 43820 7668
rect 42404 7564 42886 7658
rect 43022 7574 43820 7658
rect 43956 7588 45662 7668
rect 45774 7670 48454 7678
rect 45774 7588 46580 7670
rect 43956 7580 46580 7588
rect 46692 7594 48454 7670
rect 48560 7690 52632 7696
rect 48560 7594 49416 7690
rect 46692 7588 49416 7594
rect 49522 7684 52632 7690
rect 49522 7682 51940 7684
rect 49522 7590 50994 7682
rect 51084 7592 51940 7682
rect 52030 7592 52632 7684
rect 51084 7590 52632 7592
rect 49522 7588 52632 7590
rect 46692 7580 52632 7588
rect 43956 7574 52632 7580
rect 43022 7564 52632 7574
rect 42404 7556 52632 7564
rect 42404 7548 44526 7556
rect 47168 7552 52632 7556
rect 50162 7548 52632 7552
rect 52932 7696 63160 7708
rect 52932 7678 58982 7696
rect 52932 7668 56190 7678
rect 52932 7658 54348 7668
rect 52932 7564 53414 7658
rect 53550 7574 54348 7658
rect 54484 7588 56190 7668
rect 56302 7670 58982 7678
rect 56302 7588 57108 7670
rect 54484 7580 57108 7588
rect 57220 7594 58982 7670
rect 59088 7690 63160 7696
rect 59088 7594 59944 7690
rect 57220 7588 59944 7594
rect 60050 7684 63160 7690
rect 60050 7682 62468 7684
rect 60050 7590 61522 7682
rect 61612 7592 62468 7682
rect 62558 7592 63160 7684
rect 61612 7590 63160 7592
rect 60050 7588 63160 7590
rect 57220 7580 63160 7588
rect 54484 7574 63160 7580
rect 53550 7564 63160 7574
rect 52932 7556 63160 7564
rect 52932 7548 55054 7556
rect 57696 7552 63160 7556
rect 60690 7548 63160 7552
rect 10646 7360 10742 7394
rect 12644 7360 12740 7394
rect 10646 7298 10680 7360
rect 12706 7298 12740 7360
rect 10646 5062 10680 5124
rect 12706 5062 12740 5124
rect 10646 5028 10742 5062
rect 12644 5028 12740 5062
rect 13400 7354 13496 7388
rect 15398 7354 15494 7388
rect 13400 7292 13434 7354
rect 15460 7292 15494 7354
rect 13400 5056 13434 5118
rect 15460 5056 15494 5118
rect 13400 5022 13496 5056
rect 15398 5022 15494 5056
rect 16216 7328 16312 7362
rect 18214 7328 18310 7362
rect 16216 7266 16250 7328
rect 18276 7266 18310 7328
rect 16216 5030 16250 5092
rect 18276 5030 18310 5092
rect 16216 4996 16312 5030
rect 18214 4996 18310 5030
rect 18740 7350 18836 7384
rect 20738 7350 20834 7384
rect 18740 7288 18774 7350
rect 20800 7288 20834 7350
rect 18740 5052 18774 5114
rect 20800 5052 20834 5114
rect 18740 5018 18836 5052
rect 20738 5018 20834 5052
rect 21254 7360 21350 7394
rect 23252 7360 23348 7394
rect 21254 7298 21288 7360
rect 23314 7298 23348 7360
rect 21254 5062 21288 5124
rect 23314 5062 23348 5124
rect 21254 5028 21350 5062
rect 23252 5028 23348 5062
rect 24008 7354 24104 7388
rect 26006 7354 26102 7388
rect 24008 7292 24042 7354
rect 26068 7292 26102 7354
rect 24008 5056 24042 5118
rect 26068 5056 26102 5118
rect 24008 5022 24104 5056
rect 26006 5022 26102 5056
rect 26824 7328 26920 7362
rect 28822 7328 28918 7362
rect 26824 7266 26858 7328
rect 28884 7266 28918 7328
rect 26824 5030 26858 5092
rect 28884 5030 28918 5092
rect 26824 4996 26920 5030
rect 28822 4996 28918 5030
rect 29348 7350 29444 7384
rect 31346 7350 31442 7384
rect 29348 7288 29382 7350
rect 31408 7288 31442 7350
rect 29348 5052 29382 5114
rect 31408 5052 31442 5114
rect 29348 5018 29444 5052
rect 31346 5018 31442 5052
rect 31782 7360 31878 7394
rect 33780 7360 33876 7394
rect 31782 7298 31816 7360
rect 33842 7298 33876 7360
rect 31782 5062 31816 5124
rect 33842 5062 33876 5124
rect 31782 5028 31878 5062
rect 33780 5028 33876 5062
rect 34536 7354 34632 7388
rect 36534 7354 36630 7388
rect 34536 7292 34570 7354
rect 36596 7292 36630 7354
rect 34536 5056 34570 5118
rect 36596 5056 36630 5118
rect 34536 5022 34632 5056
rect 36534 5022 36630 5056
rect 37352 7328 37448 7362
rect 39350 7328 39446 7362
rect 37352 7266 37386 7328
rect 39412 7266 39446 7328
rect 37352 5030 37386 5092
rect 39412 5030 39446 5092
rect 37352 4996 37448 5030
rect 39350 4996 39446 5030
rect 39876 7350 39972 7384
rect 41874 7350 41970 7384
rect 39876 7288 39910 7350
rect 41936 7288 41970 7350
rect 39876 5052 39910 5114
rect 41936 5052 41970 5114
rect 39876 5018 39972 5052
rect 41874 5018 41970 5052
rect 42392 7360 42488 7394
rect 44390 7360 44486 7394
rect 42392 7298 42426 7360
rect 44452 7298 44486 7360
rect 42392 5062 42426 5124
rect 44452 5062 44486 5124
rect 42392 5028 42488 5062
rect 44390 5028 44486 5062
rect 45146 7354 45242 7388
rect 47144 7354 47240 7388
rect 45146 7292 45180 7354
rect 47206 7292 47240 7354
rect 45146 5056 45180 5118
rect 47206 5056 47240 5118
rect 45146 5022 45242 5056
rect 47144 5022 47240 5056
rect 47962 7328 48058 7362
rect 49960 7328 50056 7362
rect 47962 7266 47996 7328
rect 50022 7266 50056 7328
rect 47962 5030 47996 5092
rect 50022 5030 50056 5092
rect 47962 4996 48058 5030
rect 49960 4996 50056 5030
rect 50486 7350 50582 7384
rect 52484 7350 52580 7384
rect 50486 7288 50520 7350
rect 52546 7288 52580 7350
rect 50486 5052 50520 5114
rect 52546 5052 52580 5114
rect 50486 5018 50582 5052
rect 52484 5018 52580 5052
rect 52920 7360 53016 7394
rect 54918 7360 55014 7394
rect 52920 7298 52954 7360
rect 54980 7298 55014 7360
rect 52920 5062 52954 5124
rect 54980 5062 55014 5124
rect 52920 5028 53016 5062
rect 54918 5028 55014 5062
rect 55674 7354 55770 7388
rect 57672 7354 57768 7388
rect 55674 7292 55708 7354
rect 57734 7292 57768 7354
rect 55674 5056 55708 5118
rect 57734 5056 57768 5118
rect 55674 5022 55770 5056
rect 57672 5022 57768 5056
rect 58490 7328 58586 7362
rect 60488 7328 60584 7362
rect 58490 7266 58524 7328
rect 60550 7266 60584 7328
rect 58490 5030 58524 5092
rect 60550 5030 60584 5092
rect 58490 4996 58586 5030
rect 60488 4996 60584 5030
rect 61014 7350 61110 7384
rect 63012 7350 63108 7384
rect 61014 7288 61048 7350
rect 63074 7288 63108 7350
rect 61014 5052 61048 5114
rect 63074 5052 63108 5114
rect 61014 5018 61110 5052
rect 63012 5018 63108 5052
<< psubdiffcont >>
rect 12002 4202 14158 4236
rect 11906 3982 11940 4140
rect 14220 3982 14254 4140
rect 12002 3886 14158 3920
rect 17452 4212 19608 4246
rect 17356 3992 17390 4150
rect 19670 3992 19704 4150
rect 17452 3896 19608 3930
rect 22610 4202 24766 4236
rect 22514 3982 22548 4140
rect 24828 3982 24862 4140
rect 22610 3886 24766 3920
rect 28060 4212 30216 4246
rect 27964 3992 27998 4150
rect 30278 3992 30312 4150
rect 28060 3896 30216 3930
rect 33138 4202 35294 4236
rect 33042 3982 33076 4140
rect 35356 3982 35390 4140
rect 33138 3886 35294 3920
rect 38588 4212 40744 4246
rect 38492 3992 38526 4150
rect 40806 3992 40840 4150
rect 38588 3896 40744 3930
rect 43748 4202 45904 4236
rect 43652 3982 43686 4140
rect 45966 3982 46000 4140
rect 43748 3886 45904 3920
rect 49198 4212 51354 4246
rect 49102 3992 49136 4150
rect 51416 3992 51450 4150
rect 49198 3896 51354 3930
rect 54276 4202 56432 4236
rect 54180 3982 54214 4140
rect 56494 3982 56528 4140
rect 54276 3886 56432 3920
rect 59726 4212 61882 4246
rect 59630 3992 59664 4150
rect 61944 3992 61978 4150
rect 59726 3896 61882 3930
rect 14411 3193 19519 3227
rect 14315 575 14349 3131
rect 19581 575 19615 3131
rect 14411 479 19519 513
rect 25019 3193 30127 3227
rect 24923 575 24957 3131
rect 30189 575 30223 3131
rect 25019 479 30127 513
rect 35547 3193 40655 3227
rect 35451 575 35485 3131
rect 40717 575 40751 3131
rect 35547 479 40655 513
rect 46157 3193 51265 3227
rect 46061 575 46095 3131
rect 51327 575 51361 3131
rect 46157 479 51265 513
rect 56685 3193 61793 3227
rect 56589 575 56623 3131
rect 61855 575 61889 3131
rect 56685 479 61793 513
rect 14828 142 14986 258
rect 15722 148 15880 264
rect 17492 148 17650 264
rect 18590 152 18748 268
rect 25436 142 25594 258
rect 26330 148 26488 264
rect 28100 148 28258 264
rect 29198 152 29356 268
rect 35964 142 36122 258
rect 36858 148 37016 264
rect 38628 148 38786 264
rect 39726 152 39884 268
rect 46574 142 46732 258
rect 47468 148 47626 264
rect 49238 148 49396 264
rect 50336 152 50494 268
rect 57102 142 57260 258
rect 57996 148 58154 264
rect 59766 148 59924 264
rect 60864 152 61022 268
<< nsubdiffcont >>
rect 11140 7564 11276 7658
rect 12074 7574 12210 7668
rect 13916 7588 14028 7678
rect 14834 7580 14946 7670
rect 16708 7594 16814 7696
rect 17670 7588 17776 7690
rect 19248 7590 19338 7682
rect 20194 7592 20284 7684
rect 21748 7564 21884 7658
rect 22682 7574 22818 7668
rect 24524 7588 24636 7678
rect 25442 7580 25554 7670
rect 27316 7594 27422 7696
rect 28278 7588 28384 7690
rect 29856 7590 29946 7682
rect 30802 7592 30892 7684
rect 32276 7564 32412 7658
rect 33210 7574 33346 7668
rect 35052 7588 35164 7678
rect 35970 7580 36082 7670
rect 37844 7594 37950 7696
rect 38806 7588 38912 7690
rect 40384 7590 40474 7682
rect 41330 7592 41420 7684
rect 42886 7564 43022 7658
rect 43820 7574 43956 7668
rect 45662 7588 45774 7678
rect 46580 7580 46692 7670
rect 48454 7594 48560 7696
rect 49416 7588 49522 7690
rect 50994 7590 51084 7682
rect 51940 7592 52030 7684
rect 53414 7564 53550 7658
rect 54348 7574 54484 7668
rect 56190 7588 56302 7678
rect 57108 7580 57220 7670
rect 58982 7594 59088 7696
rect 59944 7588 60050 7690
rect 61522 7590 61612 7682
rect 62468 7592 62558 7684
rect 10742 7360 12644 7394
rect 10646 5124 10680 7298
rect 12706 5124 12740 7298
rect 10742 5028 12644 5062
rect 13496 7354 15398 7388
rect 13400 5118 13434 7292
rect 15460 5118 15494 7292
rect 13496 5022 15398 5056
rect 16312 7328 18214 7362
rect 16216 5092 16250 7266
rect 18276 5092 18310 7266
rect 16312 4996 18214 5030
rect 18836 7350 20738 7384
rect 18740 5114 18774 7288
rect 20800 5114 20834 7288
rect 18836 5018 20738 5052
rect 21350 7360 23252 7394
rect 21254 5124 21288 7298
rect 23314 5124 23348 7298
rect 21350 5028 23252 5062
rect 24104 7354 26006 7388
rect 24008 5118 24042 7292
rect 26068 5118 26102 7292
rect 24104 5022 26006 5056
rect 26920 7328 28822 7362
rect 26824 5092 26858 7266
rect 28884 5092 28918 7266
rect 26920 4996 28822 5030
rect 29444 7350 31346 7384
rect 29348 5114 29382 7288
rect 31408 5114 31442 7288
rect 29444 5018 31346 5052
rect 31878 7360 33780 7394
rect 31782 5124 31816 7298
rect 33842 5124 33876 7298
rect 31878 5028 33780 5062
rect 34632 7354 36534 7388
rect 34536 5118 34570 7292
rect 36596 5118 36630 7292
rect 34632 5022 36534 5056
rect 37448 7328 39350 7362
rect 37352 5092 37386 7266
rect 39412 5092 39446 7266
rect 37448 4996 39350 5030
rect 39972 7350 41874 7384
rect 39876 5114 39910 7288
rect 41936 5114 41970 7288
rect 39972 5018 41874 5052
rect 42488 7360 44390 7394
rect 42392 5124 42426 7298
rect 44452 5124 44486 7298
rect 42488 5028 44390 5062
rect 45242 7354 47144 7388
rect 45146 5118 45180 7292
rect 47206 5118 47240 7292
rect 45242 5022 47144 5056
rect 48058 7328 49960 7362
rect 47962 5092 47996 7266
rect 50022 5092 50056 7266
rect 48058 4996 49960 5030
rect 50582 7350 52484 7384
rect 50486 5114 50520 7288
rect 52546 5114 52580 7288
rect 50582 5018 52484 5052
rect 53016 7360 54918 7394
rect 52920 5124 52954 7298
rect 54980 5124 55014 7298
rect 53016 5028 54918 5062
rect 55770 7354 57672 7388
rect 55674 5118 55708 7292
rect 57734 5118 57768 7292
rect 55770 5022 57672 5056
rect 58586 7328 60488 7362
rect 58490 5092 58524 7266
rect 60550 5092 60584 7266
rect 58586 4996 60488 5030
rect 61110 7350 63012 7384
rect 61014 5114 61048 7288
rect 63074 5114 63108 7288
rect 61110 5018 63012 5052
<< poly >>
rect 10806 7292 11206 7308
rect 10806 7258 10822 7292
rect 11190 7258 11206 7292
rect 10806 7211 11206 7258
rect 11264 7292 11664 7308
rect 11264 7258 11280 7292
rect 11648 7258 11664 7292
rect 11264 7211 11664 7258
rect 11722 7292 12122 7308
rect 11722 7258 11738 7292
rect 12106 7258 12122 7292
rect 11722 7211 12122 7258
rect 12180 7292 12580 7308
rect 12180 7258 12196 7292
rect 12564 7258 12580 7292
rect 12180 7211 12580 7258
rect 10806 5164 11206 5211
rect 10806 5130 10822 5164
rect 11190 5130 11206 5164
rect 10806 5114 11206 5130
rect 11264 5164 11664 5211
rect 11264 5130 11280 5164
rect 11648 5130 11664 5164
rect 11264 5114 11664 5130
rect 11722 5164 12122 5211
rect 11722 5130 11738 5164
rect 12106 5130 12122 5164
rect 11722 5114 12122 5130
rect 12180 5164 12580 5211
rect 12180 5130 12196 5164
rect 12564 5130 12580 5164
rect 12180 5114 12580 5130
rect 13560 7286 13960 7302
rect 13560 7252 13576 7286
rect 13944 7252 13960 7286
rect 13560 7205 13960 7252
rect 14018 7286 14418 7302
rect 14018 7252 14034 7286
rect 14402 7252 14418 7286
rect 14018 7205 14418 7252
rect 14476 7286 14876 7302
rect 14476 7252 14492 7286
rect 14860 7252 14876 7286
rect 14476 7205 14876 7252
rect 14934 7286 15334 7302
rect 14934 7252 14950 7286
rect 15318 7252 15334 7286
rect 14934 7205 15334 7252
rect 13560 5158 13960 5205
rect 13560 5124 13576 5158
rect 13944 5124 13960 5158
rect 13560 5108 13960 5124
rect 14018 5158 14418 5205
rect 14018 5124 14034 5158
rect 14402 5124 14418 5158
rect 14018 5108 14418 5124
rect 14476 5158 14876 5205
rect 14476 5124 14492 5158
rect 14860 5124 14876 5158
rect 14476 5108 14876 5124
rect 14934 5158 15334 5205
rect 14934 5124 14950 5158
rect 15318 5124 15334 5158
rect 14934 5108 15334 5124
rect 16376 7260 16776 7276
rect 16376 7226 16392 7260
rect 16760 7226 16776 7260
rect 16376 7179 16776 7226
rect 16834 7260 17234 7276
rect 16834 7226 16850 7260
rect 17218 7226 17234 7260
rect 16834 7179 17234 7226
rect 17292 7260 17692 7276
rect 17292 7226 17308 7260
rect 17676 7226 17692 7260
rect 17292 7179 17692 7226
rect 17750 7260 18150 7276
rect 17750 7226 17766 7260
rect 18134 7226 18150 7260
rect 17750 7179 18150 7226
rect 16376 5132 16776 5179
rect 16376 5098 16392 5132
rect 16760 5098 16776 5132
rect 16376 5082 16776 5098
rect 16834 5132 17234 5179
rect 16834 5098 16850 5132
rect 17218 5098 17234 5132
rect 16834 5082 17234 5098
rect 17292 5132 17692 5179
rect 17292 5098 17308 5132
rect 17676 5098 17692 5132
rect 17292 5082 17692 5098
rect 17750 5132 18150 5179
rect 17750 5098 17766 5132
rect 18134 5098 18150 5132
rect 17750 5082 18150 5098
rect 18900 7282 19300 7298
rect 18900 7248 18916 7282
rect 19284 7248 19300 7282
rect 18900 7201 19300 7248
rect 19358 7282 19758 7298
rect 19358 7248 19374 7282
rect 19742 7248 19758 7282
rect 19358 7201 19758 7248
rect 19816 7282 20216 7298
rect 19816 7248 19832 7282
rect 20200 7248 20216 7282
rect 19816 7201 20216 7248
rect 20274 7282 20674 7298
rect 20274 7248 20290 7282
rect 20658 7248 20674 7282
rect 20274 7201 20674 7248
rect 18900 5154 19300 5201
rect 18900 5120 18916 5154
rect 19284 5120 19300 5154
rect 18900 5104 19300 5120
rect 19358 5154 19758 5201
rect 19358 5120 19374 5154
rect 19742 5120 19758 5154
rect 19358 5104 19758 5120
rect 19816 5154 20216 5201
rect 19816 5120 19832 5154
rect 20200 5120 20216 5154
rect 19816 5104 20216 5120
rect 20274 5154 20674 5201
rect 20274 5120 20290 5154
rect 20658 5120 20674 5154
rect 20274 5104 20674 5120
rect 21414 7292 21814 7308
rect 21414 7258 21430 7292
rect 21798 7258 21814 7292
rect 21414 7211 21814 7258
rect 21872 7292 22272 7308
rect 21872 7258 21888 7292
rect 22256 7258 22272 7292
rect 21872 7211 22272 7258
rect 22330 7292 22730 7308
rect 22330 7258 22346 7292
rect 22714 7258 22730 7292
rect 22330 7211 22730 7258
rect 22788 7292 23188 7308
rect 22788 7258 22804 7292
rect 23172 7258 23188 7292
rect 22788 7211 23188 7258
rect 21414 5164 21814 5211
rect 21414 5130 21430 5164
rect 21798 5130 21814 5164
rect 21414 5114 21814 5130
rect 21872 5164 22272 5211
rect 21872 5130 21888 5164
rect 22256 5130 22272 5164
rect 21872 5114 22272 5130
rect 22330 5164 22730 5211
rect 22330 5130 22346 5164
rect 22714 5130 22730 5164
rect 22330 5114 22730 5130
rect 22788 5164 23188 5211
rect 22788 5130 22804 5164
rect 23172 5130 23188 5164
rect 22788 5114 23188 5130
rect 24168 7286 24568 7302
rect 24168 7252 24184 7286
rect 24552 7252 24568 7286
rect 24168 7205 24568 7252
rect 24626 7286 25026 7302
rect 24626 7252 24642 7286
rect 25010 7252 25026 7286
rect 24626 7205 25026 7252
rect 25084 7286 25484 7302
rect 25084 7252 25100 7286
rect 25468 7252 25484 7286
rect 25084 7205 25484 7252
rect 25542 7286 25942 7302
rect 25542 7252 25558 7286
rect 25926 7252 25942 7286
rect 25542 7205 25942 7252
rect 24168 5158 24568 5205
rect 24168 5124 24184 5158
rect 24552 5124 24568 5158
rect 24168 5108 24568 5124
rect 24626 5158 25026 5205
rect 24626 5124 24642 5158
rect 25010 5124 25026 5158
rect 24626 5108 25026 5124
rect 25084 5158 25484 5205
rect 25084 5124 25100 5158
rect 25468 5124 25484 5158
rect 25084 5108 25484 5124
rect 25542 5158 25942 5205
rect 25542 5124 25558 5158
rect 25926 5124 25942 5158
rect 25542 5108 25942 5124
rect 26984 7260 27384 7276
rect 26984 7226 27000 7260
rect 27368 7226 27384 7260
rect 26984 7179 27384 7226
rect 27442 7260 27842 7276
rect 27442 7226 27458 7260
rect 27826 7226 27842 7260
rect 27442 7179 27842 7226
rect 27900 7260 28300 7276
rect 27900 7226 27916 7260
rect 28284 7226 28300 7260
rect 27900 7179 28300 7226
rect 28358 7260 28758 7276
rect 28358 7226 28374 7260
rect 28742 7226 28758 7260
rect 28358 7179 28758 7226
rect 26984 5132 27384 5179
rect 26984 5098 27000 5132
rect 27368 5098 27384 5132
rect 26984 5082 27384 5098
rect 27442 5132 27842 5179
rect 27442 5098 27458 5132
rect 27826 5098 27842 5132
rect 27442 5082 27842 5098
rect 27900 5132 28300 5179
rect 27900 5098 27916 5132
rect 28284 5098 28300 5132
rect 27900 5082 28300 5098
rect 28358 5132 28758 5179
rect 28358 5098 28374 5132
rect 28742 5098 28758 5132
rect 28358 5082 28758 5098
rect 29508 7282 29908 7298
rect 29508 7248 29524 7282
rect 29892 7248 29908 7282
rect 29508 7201 29908 7248
rect 29966 7282 30366 7298
rect 29966 7248 29982 7282
rect 30350 7248 30366 7282
rect 29966 7201 30366 7248
rect 30424 7282 30824 7298
rect 30424 7248 30440 7282
rect 30808 7248 30824 7282
rect 30424 7201 30824 7248
rect 30882 7282 31282 7298
rect 30882 7248 30898 7282
rect 31266 7248 31282 7282
rect 30882 7201 31282 7248
rect 29508 5154 29908 5201
rect 29508 5120 29524 5154
rect 29892 5120 29908 5154
rect 29508 5104 29908 5120
rect 29966 5154 30366 5201
rect 29966 5120 29982 5154
rect 30350 5120 30366 5154
rect 29966 5104 30366 5120
rect 30424 5154 30824 5201
rect 30424 5120 30440 5154
rect 30808 5120 30824 5154
rect 30424 5104 30824 5120
rect 30882 5154 31282 5201
rect 30882 5120 30898 5154
rect 31266 5120 31282 5154
rect 30882 5104 31282 5120
rect 31942 7292 32342 7308
rect 31942 7258 31958 7292
rect 32326 7258 32342 7292
rect 31942 7211 32342 7258
rect 32400 7292 32800 7308
rect 32400 7258 32416 7292
rect 32784 7258 32800 7292
rect 32400 7211 32800 7258
rect 32858 7292 33258 7308
rect 32858 7258 32874 7292
rect 33242 7258 33258 7292
rect 32858 7211 33258 7258
rect 33316 7292 33716 7308
rect 33316 7258 33332 7292
rect 33700 7258 33716 7292
rect 33316 7211 33716 7258
rect 31942 5164 32342 5211
rect 31942 5130 31958 5164
rect 32326 5130 32342 5164
rect 31942 5114 32342 5130
rect 32400 5164 32800 5211
rect 32400 5130 32416 5164
rect 32784 5130 32800 5164
rect 32400 5114 32800 5130
rect 32858 5164 33258 5211
rect 32858 5130 32874 5164
rect 33242 5130 33258 5164
rect 32858 5114 33258 5130
rect 33316 5164 33716 5211
rect 33316 5130 33332 5164
rect 33700 5130 33716 5164
rect 33316 5114 33716 5130
rect 34696 7286 35096 7302
rect 34696 7252 34712 7286
rect 35080 7252 35096 7286
rect 34696 7205 35096 7252
rect 35154 7286 35554 7302
rect 35154 7252 35170 7286
rect 35538 7252 35554 7286
rect 35154 7205 35554 7252
rect 35612 7286 36012 7302
rect 35612 7252 35628 7286
rect 35996 7252 36012 7286
rect 35612 7205 36012 7252
rect 36070 7286 36470 7302
rect 36070 7252 36086 7286
rect 36454 7252 36470 7286
rect 36070 7205 36470 7252
rect 34696 5158 35096 5205
rect 34696 5124 34712 5158
rect 35080 5124 35096 5158
rect 34696 5108 35096 5124
rect 35154 5158 35554 5205
rect 35154 5124 35170 5158
rect 35538 5124 35554 5158
rect 35154 5108 35554 5124
rect 35612 5158 36012 5205
rect 35612 5124 35628 5158
rect 35996 5124 36012 5158
rect 35612 5108 36012 5124
rect 36070 5158 36470 5205
rect 36070 5124 36086 5158
rect 36454 5124 36470 5158
rect 36070 5108 36470 5124
rect 37512 7260 37912 7276
rect 37512 7226 37528 7260
rect 37896 7226 37912 7260
rect 37512 7179 37912 7226
rect 37970 7260 38370 7276
rect 37970 7226 37986 7260
rect 38354 7226 38370 7260
rect 37970 7179 38370 7226
rect 38428 7260 38828 7276
rect 38428 7226 38444 7260
rect 38812 7226 38828 7260
rect 38428 7179 38828 7226
rect 38886 7260 39286 7276
rect 38886 7226 38902 7260
rect 39270 7226 39286 7260
rect 38886 7179 39286 7226
rect 37512 5132 37912 5179
rect 37512 5098 37528 5132
rect 37896 5098 37912 5132
rect 37512 5082 37912 5098
rect 37970 5132 38370 5179
rect 37970 5098 37986 5132
rect 38354 5098 38370 5132
rect 37970 5082 38370 5098
rect 38428 5132 38828 5179
rect 38428 5098 38444 5132
rect 38812 5098 38828 5132
rect 38428 5082 38828 5098
rect 38886 5132 39286 5179
rect 38886 5098 38902 5132
rect 39270 5098 39286 5132
rect 38886 5082 39286 5098
rect 40036 7282 40436 7298
rect 40036 7248 40052 7282
rect 40420 7248 40436 7282
rect 40036 7201 40436 7248
rect 40494 7282 40894 7298
rect 40494 7248 40510 7282
rect 40878 7248 40894 7282
rect 40494 7201 40894 7248
rect 40952 7282 41352 7298
rect 40952 7248 40968 7282
rect 41336 7248 41352 7282
rect 40952 7201 41352 7248
rect 41410 7282 41810 7298
rect 41410 7248 41426 7282
rect 41794 7248 41810 7282
rect 41410 7201 41810 7248
rect 40036 5154 40436 5201
rect 40036 5120 40052 5154
rect 40420 5120 40436 5154
rect 40036 5104 40436 5120
rect 40494 5154 40894 5201
rect 40494 5120 40510 5154
rect 40878 5120 40894 5154
rect 40494 5104 40894 5120
rect 40952 5154 41352 5201
rect 40952 5120 40968 5154
rect 41336 5120 41352 5154
rect 40952 5104 41352 5120
rect 41410 5154 41810 5201
rect 41410 5120 41426 5154
rect 41794 5120 41810 5154
rect 41410 5104 41810 5120
rect 42552 7292 42952 7308
rect 42552 7258 42568 7292
rect 42936 7258 42952 7292
rect 42552 7211 42952 7258
rect 43010 7292 43410 7308
rect 43010 7258 43026 7292
rect 43394 7258 43410 7292
rect 43010 7211 43410 7258
rect 43468 7292 43868 7308
rect 43468 7258 43484 7292
rect 43852 7258 43868 7292
rect 43468 7211 43868 7258
rect 43926 7292 44326 7308
rect 43926 7258 43942 7292
rect 44310 7258 44326 7292
rect 43926 7211 44326 7258
rect 42552 5164 42952 5211
rect 42552 5130 42568 5164
rect 42936 5130 42952 5164
rect 42552 5114 42952 5130
rect 43010 5164 43410 5211
rect 43010 5130 43026 5164
rect 43394 5130 43410 5164
rect 43010 5114 43410 5130
rect 43468 5164 43868 5211
rect 43468 5130 43484 5164
rect 43852 5130 43868 5164
rect 43468 5114 43868 5130
rect 43926 5164 44326 5211
rect 43926 5130 43942 5164
rect 44310 5130 44326 5164
rect 43926 5114 44326 5130
rect 45306 7286 45706 7302
rect 45306 7252 45322 7286
rect 45690 7252 45706 7286
rect 45306 7205 45706 7252
rect 45764 7286 46164 7302
rect 45764 7252 45780 7286
rect 46148 7252 46164 7286
rect 45764 7205 46164 7252
rect 46222 7286 46622 7302
rect 46222 7252 46238 7286
rect 46606 7252 46622 7286
rect 46222 7205 46622 7252
rect 46680 7286 47080 7302
rect 46680 7252 46696 7286
rect 47064 7252 47080 7286
rect 46680 7205 47080 7252
rect 45306 5158 45706 5205
rect 45306 5124 45322 5158
rect 45690 5124 45706 5158
rect 45306 5108 45706 5124
rect 45764 5158 46164 5205
rect 45764 5124 45780 5158
rect 46148 5124 46164 5158
rect 45764 5108 46164 5124
rect 46222 5158 46622 5205
rect 46222 5124 46238 5158
rect 46606 5124 46622 5158
rect 46222 5108 46622 5124
rect 46680 5158 47080 5205
rect 46680 5124 46696 5158
rect 47064 5124 47080 5158
rect 46680 5108 47080 5124
rect 48122 7260 48522 7276
rect 48122 7226 48138 7260
rect 48506 7226 48522 7260
rect 48122 7179 48522 7226
rect 48580 7260 48980 7276
rect 48580 7226 48596 7260
rect 48964 7226 48980 7260
rect 48580 7179 48980 7226
rect 49038 7260 49438 7276
rect 49038 7226 49054 7260
rect 49422 7226 49438 7260
rect 49038 7179 49438 7226
rect 49496 7260 49896 7276
rect 49496 7226 49512 7260
rect 49880 7226 49896 7260
rect 49496 7179 49896 7226
rect 48122 5132 48522 5179
rect 48122 5098 48138 5132
rect 48506 5098 48522 5132
rect 48122 5082 48522 5098
rect 48580 5132 48980 5179
rect 48580 5098 48596 5132
rect 48964 5098 48980 5132
rect 48580 5082 48980 5098
rect 49038 5132 49438 5179
rect 49038 5098 49054 5132
rect 49422 5098 49438 5132
rect 49038 5082 49438 5098
rect 49496 5132 49896 5179
rect 49496 5098 49512 5132
rect 49880 5098 49896 5132
rect 49496 5082 49896 5098
rect 50646 7282 51046 7298
rect 50646 7248 50662 7282
rect 51030 7248 51046 7282
rect 50646 7201 51046 7248
rect 51104 7282 51504 7298
rect 51104 7248 51120 7282
rect 51488 7248 51504 7282
rect 51104 7201 51504 7248
rect 51562 7282 51962 7298
rect 51562 7248 51578 7282
rect 51946 7248 51962 7282
rect 51562 7201 51962 7248
rect 52020 7282 52420 7298
rect 52020 7248 52036 7282
rect 52404 7248 52420 7282
rect 52020 7201 52420 7248
rect 50646 5154 51046 5201
rect 50646 5120 50662 5154
rect 51030 5120 51046 5154
rect 50646 5104 51046 5120
rect 51104 5154 51504 5201
rect 51104 5120 51120 5154
rect 51488 5120 51504 5154
rect 51104 5104 51504 5120
rect 51562 5154 51962 5201
rect 51562 5120 51578 5154
rect 51946 5120 51962 5154
rect 51562 5104 51962 5120
rect 52020 5154 52420 5201
rect 52020 5120 52036 5154
rect 52404 5120 52420 5154
rect 52020 5104 52420 5120
rect 53080 7292 53480 7308
rect 53080 7258 53096 7292
rect 53464 7258 53480 7292
rect 53080 7211 53480 7258
rect 53538 7292 53938 7308
rect 53538 7258 53554 7292
rect 53922 7258 53938 7292
rect 53538 7211 53938 7258
rect 53996 7292 54396 7308
rect 53996 7258 54012 7292
rect 54380 7258 54396 7292
rect 53996 7211 54396 7258
rect 54454 7292 54854 7308
rect 54454 7258 54470 7292
rect 54838 7258 54854 7292
rect 54454 7211 54854 7258
rect 53080 5164 53480 5211
rect 53080 5130 53096 5164
rect 53464 5130 53480 5164
rect 53080 5114 53480 5130
rect 53538 5164 53938 5211
rect 53538 5130 53554 5164
rect 53922 5130 53938 5164
rect 53538 5114 53938 5130
rect 53996 5164 54396 5211
rect 53996 5130 54012 5164
rect 54380 5130 54396 5164
rect 53996 5114 54396 5130
rect 54454 5164 54854 5211
rect 54454 5130 54470 5164
rect 54838 5130 54854 5164
rect 54454 5114 54854 5130
rect 55834 7286 56234 7302
rect 55834 7252 55850 7286
rect 56218 7252 56234 7286
rect 55834 7205 56234 7252
rect 56292 7286 56692 7302
rect 56292 7252 56308 7286
rect 56676 7252 56692 7286
rect 56292 7205 56692 7252
rect 56750 7286 57150 7302
rect 56750 7252 56766 7286
rect 57134 7252 57150 7286
rect 56750 7205 57150 7252
rect 57208 7286 57608 7302
rect 57208 7252 57224 7286
rect 57592 7252 57608 7286
rect 57208 7205 57608 7252
rect 55834 5158 56234 5205
rect 55834 5124 55850 5158
rect 56218 5124 56234 5158
rect 55834 5108 56234 5124
rect 56292 5158 56692 5205
rect 56292 5124 56308 5158
rect 56676 5124 56692 5158
rect 56292 5108 56692 5124
rect 56750 5158 57150 5205
rect 56750 5124 56766 5158
rect 57134 5124 57150 5158
rect 56750 5108 57150 5124
rect 57208 5158 57608 5205
rect 57208 5124 57224 5158
rect 57592 5124 57608 5158
rect 57208 5108 57608 5124
rect 58650 7260 59050 7276
rect 58650 7226 58666 7260
rect 59034 7226 59050 7260
rect 58650 7179 59050 7226
rect 59108 7260 59508 7276
rect 59108 7226 59124 7260
rect 59492 7226 59508 7260
rect 59108 7179 59508 7226
rect 59566 7260 59966 7276
rect 59566 7226 59582 7260
rect 59950 7226 59966 7260
rect 59566 7179 59966 7226
rect 60024 7260 60424 7276
rect 60024 7226 60040 7260
rect 60408 7226 60424 7260
rect 60024 7179 60424 7226
rect 58650 5132 59050 5179
rect 58650 5098 58666 5132
rect 59034 5098 59050 5132
rect 58650 5082 59050 5098
rect 59108 5132 59508 5179
rect 59108 5098 59124 5132
rect 59492 5098 59508 5132
rect 59108 5082 59508 5098
rect 59566 5132 59966 5179
rect 59566 5098 59582 5132
rect 59950 5098 59966 5132
rect 59566 5082 59966 5098
rect 60024 5132 60424 5179
rect 60024 5098 60040 5132
rect 60408 5098 60424 5132
rect 60024 5082 60424 5098
rect 61174 7282 61574 7298
rect 61174 7248 61190 7282
rect 61558 7248 61574 7282
rect 61174 7201 61574 7248
rect 61632 7282 62032 7298
rect 61632 7248 61648 7282
rect 62016 7248 62032 7282
rect 61632 7201 62032 7248
rect 62090 7282 62490 7298
rect 62090 7248 62106 7282
rect 62474 7248 62490 7282
rect 62090 7201 62490 7248
rect 62548 7282 62948 7298
rect 62548 7248 62564 7282
rect 62932 7248 62948 7282
rect 62548 7201 62948 7248
rect 61174 5154 61574 5201
rect 61174 5120 61190 5154
rect 61558 5120 61574 5154
rect 61174 5104 61574 5120
rect 61632 5154 62032 5201
rect 61632 5120 61648 5154
rect 62016 5120 62032 5154
rect 61632 5104 62032 5120
rect 62090 5154 62490 5201
rect 62090 5120 62106 5154
rect 62474 5120 62490 5154
rect 62090 5104 62490 5120
rect 62548 5154 62948 5201
rect 62548 5120 62564 5154
rect 62932 5120 62948 5154
rect 62548 5104 62948 5120
rect 11992 4078 12058 4094
rect 11992 4044 12008 4078
rect 12042 4076 12058 4078
rect 14102 4078 14168 4094
rect 14102 4076 14118 4078
rect 12042 4046 12080 4076
rect 14080 4046 14118 4076
rect 12042 4044 12058 4046
rect 11992 4028 12058 4044
rect 14102 4044 14118 4046
rect 14152 4044 14168 4078
rect 14102 4028 14168 4044
rect 17442 4088 17508 4104
rect 17442 4054 17458 4088
rect 17492 4086 17508 4088
rect 19552 4088 19618 4104
rect 19552 4086 19568 4088
rect 17492 4056 17530 4086
rect 19530 4056 19568 4086
rect 17492 4054 17508 4056
rect 17442 4038 17508 4054
rect 19552 4054 19568 4056
rect 19602 4054 19618 4088
rect 19552 4038 19618 4054
rect 22600 4078 22666 4094
rect 22600 4044 22616 4078
rect 22650 4076 22666 4078
rect 24710 4078 24776 4094
rect 24710 4076 24726 4078
rect 22650 4046 22688 4076
rect 24688 4046 24726 4076
rect 22650 4044 22666 4046
rect 22600 4028 22666 4044
rect 24710 4044 24726 4046
rect 24760 4044 24776 4078
rect 24710 4028 24776 4044
rect 28050 4088 28116 4104
rect 28050 4054 28066 4088
rect 28100 4086 28116 4088
rect 30160 4088 30226 4104
rect 30160 4086 30176 4088
rect 28100 4056 28138 4086
rect 30138 4056 30176 4086
rect 28100 4054 28116 4056
rect 28050 4038 28116 4054
rect 30160 4054 30176 4056
rect 30210 4054 30226 4088
rect 30160 4038 30226 4054
rect 33128 4078 33194 4094
rect 33128 4044 33144 4078
rect 33178 4076 33194 4078
rect 35238 4078 35304 4094
rect 35238 4076 35254 4078
rect 33178 4046 33216 4076
rect 35216 4046 35254 4076
rect 33178 4044 33194 4046
rect 33128 4028 33194 4044
rect 35238 4044 35254 4046
rect 35288 4044 35304 4078
rect 35238 4028 35304 4044
rect 38578 4088 38644 4104
rect 38578 4054 38594 4088
rect 38628 4086 38644 4088
rect 40688 4088 40754 4104
rect 40688 4086 40704 4088
rect 38628 4056 38666 4086
rect 40666 4056 40704 4086
rect 38628 4054 38644 4056
rect 38578 4038 38644 4054
rect 40688 4054 40704 4056
rect 40738 4054 40754 4088
rect 40688 4038 40754 4054
rect 43738 4078 43804 4094
rect 43738 4044 43754 4078
rect 43788 4076 43804 4078
rect 45848 4078 45914 4094
rect 45848 4076 45864 4078
rect 43788 4046 43826 4076
rect 45826 4046 45864 4076
rect 43788 4044 43804 4046
rect 43738 4028 43804 4044
rect 45848 4044 45864 4046
rect 45898 4044 45914 4078
rect 45848 4028 45914 4044
rect 49188 4088 49254 4104
rect 49188 4054 49204 4088
rect 49238 4086 49254 4088
rect 51298 4088 51364 4104
rect 51298 4086 51314 4088
rect 49238 4056 49276 4086
rect 51276 4056 51314 4086
rect 49238 4054 49254 4056
rect 49188 4038 49254 4054
rect 51298 4054 51314 4056
rect 51348 4054 51364 4088
rect 51298 4038 51364 4054
rect 54266 4078 54332 4094
rect 54266 4044 54282 4078
rect 54316 4076 54332 4078
rect 56376 4078 56442 4094
rect 56376 4076 56392 4078
rect 54316 4046 54354 4076
rect 56354 4046 56392 4076
rect 54316 4044 54332 4046
rect 54266 4028 54332 4044
rect 56376 4044 56392 4046
rect 56426 4044 56442 4078
rect 56376 4028 56442 4044
rect 59716 4088 59782 4104
rect 59716 4054 59732 4088
rect 59766 4086 59782 4088
rect 61826 4088 61892 4104
rect 61826 4086 61842 4088
rect 59766 4056 59804 4086
rect 61804 4056 61842 4086
rect 59766 4054 59782 4056
rect 59716 4038 59782 4054
rect 61826 4054 61842 4056
rect 61876 4054 61892 4088
rect 61826 4038 61892 4054
rect 14475 3125 14875 3141
rect 14475 3091 14491 3125
rect 14859 3091 14875 3125
rect 14475 3053 14875 3091
rect 14933 3125 15333 3141
rect 14933 3091 14949 3125
rect 15317 3091 15333 3125
rect 14933 3053 15333 3091
rect 15391 3125 15791 3141
rect 15391 3091 15407 3125
rect 15775 3091 15791 3125
rect 15391 3053 15791 3091
rect 15849 3125 16249 3141
rect 15849 3091 15865 3125
rect 16233 3091 16249 3125
rect 15849 3053 16249 3091
rect 16307 3125 16707 3141
rect 16307 3091 16323 3125
rect 16691 3091 16707 3125
rect 16307 3053 16707 3091
rect 16765 3125 17165 3141
rect 16765 3091 16781 3125
rect 17149 3091 17165 3125
rect 16765 3053 17165 3091
rect 17223 3125 17623 3141
rect 17223 3091 17239 3125
rect 17607 3091 17623 3125
rect 17223 3053 17623 3091
rect 17681 3125 18081 3141
rect 17681 3091 17697 3125
rect 18065 3091 18081 3125
rect 17681 3053 18081 3091
rect 18139 3125 18539 3141
rect 18139 3091 18155 3125
rect 18523 3091 18539 3125
rect 18139 3053 18539 3091
rect 18597 3125 18997 3141
rect 18597 3091 18613 3125
rect 18981 3091 18997 3125
rect 18597 3053 18997 3091
rect 19055 3125 19455 3141
rect 19055 3091 19071 3125
rect 19439 3091 19455 3125
rect 19055 3053 19455 3091
rect 14475 615 14875 653
rect 14475 581 14491 615
rect 14859 581 14875 615
rect 14475 565 14875 581
rect 14933 615 15333 653
rect 14933 581 14949 615
rect 15317 581 15333 615
rect 14933 565 15333 581
rect 15391 615 15791 653
rect 15391 581 15407 615
rect 15775 581 15791 615
rect 15391 565 15791 581
rect 15849 615 16249 653
rect 15849 581 15865 615
rect 16233 581 16249 615
rect 15849 565 16249 581
rect 16307 615 16707 653
rect 16307 581 16323 615
rect 16691 581 16707 615
rect 16307 565 16707 581
rect 16765 615 17165 653
rect 16765 581 16781 615
rect 17149 581 17165 615
rect 16765 565 17165 581
rect 17223 615 17623 653
rect 17223 581 17239 615
rect 17607 581 17623 615
rect 17223 565 17623 581
rect 17681 615 18081 653
rect 17681 581 17697 615
rect 18065 581 18081 615
rect 17681 565 18081 581
rect 18139 615 18539 653
rect 18139 581 18155 615
rect 18523 581 18539 615
rect 18139 565 18539 581
rect 18597 615 18997 653
rect 18597 581 18613 615
rect 18981 581 18997 615
rect 18597 565 18997 581
rect 19055 615 19455 653
rect 19055 581 19071 615
rect 19439 581 19455 615
rect 19055 565 19455 581
rect 25083 3125 25483 3141
rect 25083 3091 25099 3125
rect 25467 3091 25483 3125
rect 25083 3053 25483 3091
rect 25541 3125 25941 3141
rect 25541 3091 25557 3125
rect 25925 3091 25941 3125
rect 25541 3053 25941 3091
rect 25999 3125 26399 3141
rect 25999 3091 26015 3125
rect 26383 3091 26399 3125
rect 25999 3053 26399 3091
rect 26457 3125 26857 3141
rect 26457 3091 26473 3125
rect 26841 3091 26857 3125
rect 26457 3053 26857 3091
rect 26915 3125 27315 3141
rect 26915 3091 26931 3125
rect 27299 3091 27315 3125
rect 26915 3053 27315 3091
rect 27373 3125 27773 3141
rect 27373 3091 27389 3125
rect 27757 3091 27773 3125
rect 27373 3053 27773 3091
rect 27831 3125 28231 3141
rect 27831 3091 27847 3125
rect 28215 3091 28231 3125
rect 27831 3053 28231 3091
rect 28289 3125 28689 3141
rect 28289 3091 28305 3125
rect 28673 3091 28689 3125
rect 28289 3053 28689 3091
rect 28747 3125 29147 3141
rect 28747 3091 28763 3125
rect 29131 3091 29147 3125
rect 28747 3053 29147 3091
rect 29205 3125 29605 3141
rect 29205 3091 29221 3125
rect 29589 3091 29605 3125
rect 29205 3053 29605 3091
rect 29663 3125 30063 3141
rect 29663 3091 29679 3125
rect 30047 3091 30063 3125
rect 29663 3053 30063 3091
rect 25083 615 25483 653
rect 25083 581 25099 615
rect 25467 581 25483 615
rect 25083 565 25483 581
rect 25541 615 25941 653
rect 25541 581 25557 615
rect 25925 581 25941 615
rect 25541 565 25941 581
rect 25999 615 26399 653
rect 25999 581 26015 615
rect 26383 581 26399 615
rect 25999 565 26399 581
rect 26457 615 26857 653
rect 26457 581 26473 615
rect 26841 581 26857 615
rect 26457 565 26857 581
rect 26915 615 27315 653
rect 26915 581 26931 615
rect 27299 581 27315 615
rect 26915 565 27315 581
rect 27373 615 27773 653
rect 27373 581 27389 615
rect 27757 581 27773 615
rect 27373 565 27773 581
rect 27831 615 28231 653
rect 27831 581 27847 615
rect 28215 581 28231 615
rect 27831 565 28231 581
rect 28289 615 28689 653
rect 28289 581 28305 615
rect 28673 581 28689 615
rect 28289 565 28689 581
rect 28747 615 29147 653
rect 28747 581 28763 615
rect 29131 581 29147 615
rect 28747 565 29147 581
rect 29205 615 29605 653
rect 29205 581 29221 615
rect 29589 581 29605 615
rect 29205 565 29605 581
rect 29663 615 30063 653
rect 29663 581 29679 615
rect 30047 581 30063 615
rect 29663 565 30063 581
rect 35611 3125 36011 3141
rect 35611 3091 35627 3125
rect 35995 3091 36011 3125
rect 35611 3053 36011 3091
rect 36069 3125 36469 3141
rect 36069 3091 36085 3125
rect 36453 3091 36469 3125
rect 36069 3053 36469 3091
rect 36527 3125 36927 3141
rect 36527 3091 36543 3125
rect 36911 3091 36927 3125
rect 36527 3053 36927 3091
rect 36985 3125 37385 3141
rect 36985 3091 37001 3125
rect 37369 3091 37385 3125
rect 36985 3053 37385 3091
rect 37443 3125 37843 3141
rect 37443 3091 37459 3125
rect 37827 3091 37843 3125
rect 37443 3053 37843 3091
rect 37901 3125 38301 3141
rect 37901 3091 37917 3125
rect 38285 3091 38301 3125
rect 37901 3053 38301 3091
rect 38359 3125 38759 3141
rect 38359 3091 38375 3125
rect 38743 3091 38759 3125
rect 38359 3053 38759 3091
rect 38817 3125 39217 3141
rect 38817 3091 38833 3125
rect 39201 3091 39217 3125
rect 38817 3053 39217 3091
rect 39275 3125 39675 3141
rect 39275 3091 39291 3125
rect 39659 3091 39675 3125
rect 39275 3053 39675 3091
rect 39733 3125 40133 3141
rect 39733 3091 39749 3125
rect 40117 3091 40133 3125
rect 39733 3053 40133 3091
rect 40191 3125 40591 3141
rect 40191 3091 40207 3125
rect 40575 3091 40591 3125
rect 40191 3053 40591 3091
rect 35611 615 36011 653
rect 35611 581 35627 615
rect 35995 581 36011 615
rect 35611 565 36011 581
rect 36069 615 36469 653
rect 36069 581 36085 615
rect 36453 581 36469 615
rect 36069 565 36469 581
rect 36527 615 36927 653
rect 36527 581 36543 615
rect 36911 581 36927 615
rect 36527 565 36927 581
rect 36985 615 37385 653
rect 36985 581 37001 615
rect 37369 581 37385 615
rect 36985 565 37385 581
rect 37443 615 37843 653
rect 37443 581 37459 615
rect 37827 581 37843 615
rect 37443 565 37843 581
rect 37901 615 38301 653
rect 37901 581 37917 615
rect 38285 581 38301 615
rect 37901 565 38301 581
rect 38359 615 38759 653
rect 38359 581 38375 615
rect 38743 581 38759 615
rect 38359 565 38759 581
rect 38817 615 39217 653
rect 38817 581 38833 615
rect 39201 581 39217 615
rect 38817 565 39217 581
rect 39275 615 39675 653
rect 39275 581 39291 615
rect 39659 581 39675 615
rect 39275 565 39675 581
rect 39733 615 40133 653
rect 39733 581 39749 615
rect 40117 581 40133 615
rect 39733 565 40133 581
rect 40191 615 40591 653
rect 40191 581 40207 615
rect 40575 581 40591 615
rect 40191 565 40591 581
rect 46221 3125 46621 3141
rect 46221 3091 46237 3125
rect 46605 3091 46621 3125
rect 46221 3053 46621 3091
rect 46679 3125 47079 3141
rect 46679 3091 46695 3125
rect 47063 3091 47079 3125
rect 46679 3053 47079 3091
rect 47137 3125 47537 3141
rect 47137 3091 47153 3125
rect 47521 3091 47537 3125
rect 47137 3053 47537 3091
rect 47595 3125 47995 3141
rect 47595 3091 47611 3125
rect 47979 3091 47995 3125
rect 47595 3053 47995 3091
rect 48053 3125 48453 3141
rect 48053 3091 48069 3125
rect 48437 3091 48453 3125
rect 48053 3053 48453 3091
rect 48511 3125 48911 3141
rect 48511 3091 48527 3125
rect 48895 3091 48911 3125
rect 48511 3053 48911 3091
rect 48969 3125 49369 3141
rect 48969 3091 48985 3125
rect 49353 3091 49369 3125
rect 48969 3053 49369 3091
rect 49427 3125 49827 3141
rect 49427 3091 49443 3125
rect 49811 3091 49827 3125
rect 49427 3053 49827 3091
rect 49885 3125 50285 3141
rect 49885 3091 49901 3125
rect 50269 3091 50285 3125
rect 49885 3053 50285 3091
rect 50343 3125 50743 3141
rect 50343 3091 50359 3125
rect 50727 3091 50743 3125
rect 50343 3053 50743 3091
rect 50801 3125 51201 3141
rect 50801 3091 50817 3125
rect 51185 3091 51201 3125
rect 50801 3053 51201 3091
rect 46221 615 46621 653
rect 46221 581 46237 615
rect 46605 581 46621 615
rect 46221 565 46621 581
rect 46679 615 47079 653
rect 46679 581 46695 615
rect 47063 581 47079 615
rect 46679 565 47079 581
rect 47137 615 47537 653
rect 47137 581 47153 615
rect 47521 581 47537 615
rect 47137 565 47537 581
rect 47595 615 47995 653
rect 47595 581 47611 615
rect 47979 581 47995 615
rect 47595 565 47995 581
rect 48053 615 48453 653
rect 48053 581 48069 615
rect 48437 581 48453 615
rect 48053 565 48453 581
rect 48511 615 48911 653
rect 48511 581 48527 615
rect 48895 581 48911 615
rect 48511 565 48911 581
rect 48969 615 49369 653
rect 48969 581 48985 615
rect 49353 581 49369 615
rect 48969 565 49369 581
rect 49427 615 49827 653
rect 49427 581 49443 615
rect 49811 581 49827 615
rect 49427 565 49827 581
rect 49885 615 50285 653
rect 49885 581 49901 615
rect 50269 581 50285 615
rect 49885 565 50285 581
rect 50343 615 50743 653
rect 50343 581 50359 615
rect 50727 581 50743 615
rect 50343 565 50743 581
rect 50801 615 51201 653
rect 50801 581 50817 615
rect 51185 581 51201 615
rect 50801 565 51201 581
rect 56749 3125 57149 3141
rect 56749 3091 56765 3125
rect 57133 3091 57149 3125
rect 56749 3053 57149 3091
rect 57207 3125 57607 3141
rect 57207 3091 57223 3125
rect 57591 3091 57607 3125
rect 57207 3053 57607 3091
rect 57665 3125 58065 3141
rect 57665 3091 57681 3125
rect 58049 3091 58065 3125
rect 57665 3053 58065 3091
rect 58123 3125 58523 3141
rect 58123 3091 58139 3125
rect 58507 3091 58523 3125
rect 58123 3053 58523 3091
rect 58581 3125 58981 3141
rect 58581 3091 58597 3125
rect 58965 3091 58981 3125
rect 58581 3053 58981 3091
rect 59039 3125 59439 3141
rect 59039 3091 59055 3125
rect 59423 3091 59439 3125
rect 59039 3053 59439 3091
rect 59497 3125 59897 3141
rect 59497 3091 59513 3125
rect 59881 3091 59897 3125
rect 59497 3053 59897 3091
rect 59955 3125 60355 3141
rect 59955 3091 59971 3125
rect 60339 3091 60355 3125
rect 59955 3053 60355 3091
rect 60413 3125 60813 3141
rect 60413 3091 60429 3125
rect 60797 3091 60813 3125
rect 60413 3053 60813 3091
rect 60871 3125 61271 3141
rect 60871 3091 60887 3125
rect 61255 3091 61271 3125
rect 60871 3053 61271 3091
rect 61329 3125 61729 3141
rect 61329 3091 61345 3125
rect 61713 3091 61729 3125
rect 61329 3053 61729 3091
rect 56749 615 57149 653
rect 56749 581 56765 615
rect 57133 581 57149 615
rect 56749 565 57149 581
rect 57207 615 57607 653
rect 57207 581 57223 615
rect 57591 581 57607 615
rect 57207 565 57607 581
rect 57665 615 58065 653
rect 57665 581 57681 615
rect 58049 581 58065 615
rect 57665 565 58065 581
rect 58123 615 58523 653
rect 58123 581 58139 615
rect 58507 581 58523 615
rect 58123 565 58523 581
rect 58581 615 58981 653
rect 58581 581 58597 615
rect 58965 581 58981 615
rect 58581 565 58981 581
rect 59039 615 59439 653
rect 59039 581 59055 615
rect 59423 581 59439 615
rect 59039 565 59439 581
rect 59497 615 59897 653
rect 59497 581 59513 615
rect 59881 581 59897 615
rect 59497 565 59897 581
rect 59955 615 60355 653
rect 59955 581 59971 615
rect 60339 581 60355 615
rect 59955 565 60355 581
rect 60413 615 60813 653
rect 60413 581 60429 615
rect 60797 581 60813 615
rect 60413 565 60813 581
rect 60871 615 61271 653
rect 60871 581 60887 615
rect 61255 581 61271 615
rect 60871 565 61271 581
rect 61329 615 61729 653
rect 61329 581 61345 615
rect 61713 581 61729 615
rect 61329 565 61729 581
<< polycont >>
rect 10822 7258 11190 7292
rect 11280 7258 11648 7292
rect 11738 7258 12106 7292
rect 12196 7258 12564 7292
rect 10822 5130 11190 5164
rect 11280 5130 11648 5164
rect 11738 5130 12106 5164
rect 12196 5130 12564 5164
rect 13576 7252 13944 7286
rect 14034 7252 14402 7286
rect 14492 7252 14860 7286
rect 14950 7252 15318 7286
rect 13576 5124 13944 5158
rect 14034 5124 14402 5158
rect 14492 5124 14860 5158
rect 14950 5124 15318 5158
rect 16392 7226 16760 7260
rect 16850 7226 17218 7260
rect 17308 7226 17676 7260
rect 17766 7226 18134 7260
rect 16392 5098 16760 5132
rect 16850 5098 17218 5132
rect 17308 5098 17676 5132
rect 17766 5098 18134 5132
rect 18916 7248 19284 7282
rect 19374 7248 19742 7282
rect 19832 7248 20200 7282
rect 20290 7248 20658 7282
rect 18916 5120 19284 5154
rect 19374 5120 19742 5154
rect 19832 5120 20200 5154
rect 20290 5120 20658 5154
rect 21430 7258 21798 7292
rect 21888 7258 22256 7292
rect 22346 7258 22714 7292
rect 22804 7258 23172 7292
rect 21430 5130 21798 5164
rect 21888 5130 22256 5164
rect 22346 5130 22714 5164
rect 22804 5130 23172 5164
rect 24184 7252 24552 7286
rect 24642 7252 25010 7286
rect 25100 7252 25468 7286
rect 25558 7252 25926 7286
rect 24184 5124 24552 5158
rect 24642 5124 25010 5158
rect 25100 5124 25468 5158
rect 25558 5124 25926 5158
rect 27000 7226 27368 7260
rect 27458 7226 27826 7260
rect 27916 7226 28284 7260
rect 28374 7226 28742 7260
rect 27000 5098 27368 5132
rect 27458 5098 27826 5132
rect 27916 5098 28284 5132
rect 28374 5098 28742 5132
rect 29524 7248 29892 7282
rect 29982 7248 30350 7282
rect 30440 7248 30808 7282
rect 30898 7248 31266 7282
rect 29524 5120 29892 5154
rect 29982 5120 30350 5154
rect 30440 5120 30808 5154
rect 30898 5120 31266 5154
rect 31958 7258 32326 7292
rect 32416 7258 32784 7292
rect 32874 7258 33242 7292
rect 33332 7258 33700 7292
rect 31958 5130 32326 5164
rect 32416 5130 32784 5164
rect 32874 5130 33242 5164
rect 33332 5130 33700 5164
rect 34712 7252 35080 7286
rect 35170 7252 35538 7286
rect 35628 7252 35996 7286
rect 36086 7252 36454 7286
rect 34712 5124 35080 5158
rect 35170 5124 35538 5158
rect 35628 5124 35996 5158
rect 36086 5124 36454 5158
rect 37528 7226 37896 7260
rect 37986 7226 38354 7260
rect 38444 7226 38812 7260
rect 38902 7226 39270 7260
rect 37528 5098 37896 5132
rect 37986 5098 38354 5132
rect 38444 5098 38812 5132
rect 38902 5098 39270 5132
rect 40052 7248 40420 7282
rect 40510 7248 40878 7282
rect 40968 7248 41336 7282
rect 41426 7248 41794 7282
rect 40052 5120 40420 5154
rect 40510 5120 40878 5154
rect 40968 5120 41336 5154
rect 41426 5120 41794 5154
rect 42568 7258 42936 7292
rect 43026 7258 43394 7292
rect 43484 7258 43852 7292
rect 43942 7258 44310 7292
rect 42568 5130 42936 5164
rect 43026 5130 43394 5164
rect 43484 5130 43852 5164
rect 43942 5130 44310 5164
rect 45322 7252 45690 7286
rect 45780 7252 46148 7286
rect 46238 7252 46606 7286
rect 46696 7252 47064 7286
rect 45322 5124 45690 5158
rect 45780 5124 46148 5158
rect 46238 5124 46606 5158
rect 46696 5124 47064 5158
rect 48138 7226 48506 7260
rect 48596 7226 48964 7260
rect 49054 7226 49422 7260
rect 49512 7226 49880 7260
rect 48138 5098 48506 5132
rect 48596 5098 48964 5132
rect 49054 5098 49422 5132
rect 49512 5098 49880 5132
rect 50662 7248 51030 7282
rect 51120 7248 51488 7282
rect 51578 7248 51946 7282
rect 52036 7248 52404 7282
rect 50662 5120 51030 5154
rect 51120 5120 51488 5154
rect 51578 5120 51946 5154
rect 52036 5120 52404 5154
rect 53096 7258 53464 7292
rect 53554 7258 53922 7292
rect 54012 7258 54380 7292
rect 54470 7258 54838 7292
rect 53096 5130 53464 5164
rect 53554 5130 53922 5164
rect 54012 5130 54380 5164
rect 54470 5130 54838 5164
rect 55850 7252 56218 7286
rect 56308 7252 56676 7286
rect 56766 7252 57134 7286
rect 57224 7252 57592 7286
rect 55850 5124 56218 5158
rect 56308 5124 56676 5158
rect 56766 5124 57134 5158
rect 57224 5124 57592 5158
rect 58666 7226 59034 7260
rect 59124 7226 59492 7260
rect 59582 7226 59950 7260
rect 60040 7226 60408 7260
rect 58666 5098 59034 5132
rect 59124 5098 59492 5132
rect 59582 5098 59950 5132
rect 60040 5098 60408 5132
rect 61190 7248 61558 7282
rect 61648 7248 62016 7282
rect 62106 7248 62474 7282
rect 62564 7248 62932 7282
rect 61190 5120 61558 5154
rect 61648 5120 62016 5154
rect 62106 5120 62474 5154
rect 62564 5120 62932 5154
rect 12008 4044 12042 4078
rect 14118 4044 14152 4078
rect 17458 4054 17492 4088
rect 19568 4054 19602 4088
rect 22616 4044 22650 4078
rect 24726 4044 24760 4078
rect 28066 4054 28100 4088
rect 30176 4054 30210 4088
rect 33144 4044 33178 4078
rect 35254 4044 35288 4078
rect 38594 4054 38628 4088
rect 40704 4054 40738 4088
rect 43754 4044 43788 4078
rect 45864 4044 45898 4078
rect 49204 4054 49238 4088
rect 51314 4054 51348 4088
rect 54282 4044 54316 4078
rect 56392 4044 56426 4078
rect 59732 4054 59766 4088
rect 61842 4054 61876 4088
rect 14491 3091 14859 3125
rect 14949 3091 15317 3125
rect 15407 3091 15775 3125
rect 15865 3091 16233 3125
rect 16323 3091 16691 3125
rect 16781 3091 17149 3125
rect 17239 3091 17607 3125
rect 17697 3091 18065 3125
rect 18155 3091 18523 3125
rect 18613 3091 18981 3125
rect 19071 3091 19439 3125
rect 14491 581 14859 615
rect 14949 581 15317 615
rect 15407 581 15775 615
rect 15865 581 16233 615
rect 16323 581 16691 615
rect 16781 581 17149 615
rect 17239 581 17607 615
rect 17697 581 18065 615
rect 18155 581 18523 615
rect 18613 581 18981 615
rect 19071 581 19439 615
rect 25099 3091 25467 3125
rect 25557 3091 25925 3125
rect 26015 3091 26383 3125
rect 26473 3091 26841 3125
rect 26931 3091 27299 3125
rect 27389 3091 27757 3125
rect 27847 3091 28215 3125
rect 28305 3091 28673 3125
rect 28763 3091 29131 3125
rect 29221 3091 29589 3125
rect 29679 3091 30047 3125
rect 25099 581 25467 615
rect 25557 581 25925 615
rect 26015 581 26383 615
rect 26473 581 26841 615
rect 26931 581 27299 615
rect 27389 581 27757 615
rect 27847 581 28215 615
rect 28305 581 28673 615
rect 28763 581 29131 615
rect 29221 581 29589 615
rect 29679 581 30047 615
rect 35627 3091 35995 3125
rect 36085 3091 36453 3125
rect 36543 3091 36911 3125
rect 37001 3091 37369 3125
rect 37459 3091 37827 3125
rect 37917 3091 38285 3125
rect 38375 3091 38743 3125
rect 38833 3091 39201 3125
rect 39291 3091 39659 3125
rect 39749 3091 40117 3125
rect 40207 3091 40575 3125
rect 35627 581 35995 615
rect 36085 581 36453 615
rect 36543 581 36911 615
rect 37001 581 37369 615
rect 37459 581 37827 615
rect 37917 581 38285 615
rect 38375 581 38743 615
rect 38833 581 39201 615
rect 39291 581 39659 615
rect 39749 581 40117 615
rect 40207 581 40575 615
rect 46237 3091 46605 3125
rect 46695 3091 47063 3125
rect 47153 3091 47521 3125
rect 47611 3091 47979 3125
rect 48069 3091 48437 3125
rect 48527 3091 48895 3125
rect 48985 3091 49353 3125
rect 49443 3091 49811 3125
rect 49901 3091 50269 3125
rect 50359 3091 50727 3125
rect 50817 3091 51185 3125
rect 46237 581 46605 615
rect 46695 581 47063 615
rect 47153 581 47521 615
rect 47611 581 47979 615
rect 48069 581 48437 615
rect 48527 581 48895 615
rect 48985 581 49353 615
rect 49443 581 49811 615
rect 49901 581 50269 615
rect 50359 581 50727 615
rect 50817 581 51185 615
rect 56765 3091 57133 3125
rect 57223 3091 57591 3125
rect 57681 3091 58049 3125
rect 58139 3091 58507 3125
rect 58597 3091 58965 3125
rect 59055 3091 59423 3125
rect 59513 3091 59881 3125
rect 59971 3091 60339 3125
rect 60429 3091 60797 3125
rect 60887 3091 61255 3125
rect 61345 3091 61713 3125
rect 56765 581 57133 615
rect 57223 581 57591 615
rect 57681 581 58049 615
rect 58139 581 58507 615
rect 58597 581 58965 615
rect 59055 581 59423 615
rect 59513 581 59881 615
rect 59971 581 60339 615
rect 60429 581 60797 615
rect 60887 581 61255 615
rect 61345 581 61713 615
<< locali >>
rect 19316 7704 20870 7708
rect 29924 7704 31478 7708
rect 40452 7704 42006 7708
rect 51062 7704 52616 7708
rect 61590 7704 63144 7708
rect 15382 7696 19740 7704
rect 15382 7688 16708 7696
rect 12674 7686 16708 7688
rect 12674 7684 16314 7686
rect 10662 7680 16314 7684
rect 10662 7678 14388 7680
rect 10662 7670 13916 7678
rect 10662 7668 13496 7670
rect 10662 7658 12074 7668
rect 10662 7646 11140 7658
rect 10662 7574 10798 7646
rect 10898 7574 11140 7646
rect 10662 7564 11140 7574
rect 11276 7654 12074 7658
rect 11276 7582 11634 7654
rect 11734 7582 12074 7654
rect 11276 7574 12074 7582
rect 12210 7666 13496 7668
rect 12210 7594 12544 7666
rect 12644 7594 13496 7666
rect 12210 7580 13496 7594
rect 13608 7588 13916 7670
rect 14028 7590 14388 7678
rect 14500 7670 16314 7680
rect 14500 7590 14834 7670
rect 14028 7588 14834 7590
rect 13608 7580 14834 7588
rect 14946 7668 16314 7670
rect 14946 7580 15278 7668
rect 12210 7578 15278 7580
rect 15390 7584 16314 7668
rect 16420 7594 16708 7686
rect 16814 7690 18828 7696
rect 16814 7676 17670 7690
rect 16814 7594 17168 7676
rect 16420 7584 17168 7594
rect 15390 7578 17168 7584
rect 12210 7576 17168 7578
rect 12210 7574 15412 7576
rect 17274 7588 17670 7676
rect 17776 7676 18828 7690
rect 17776 7588 18128 7676
rect 17274 7576 18128 7588
rect 18234 7580 18828 7676
rect 18924 7682 19740 7696
rect 18924 7590 19248 7682
rect 19338 7590 19740 7682
rect 18924 7588 19740 7590
rect 19836 7702 20870 7704
rect 19836 7684 20668 7702
rect 19836 7592 20194 7684
rect 20284 7592 20668 7684
rect 19836 7588 20668 7592
rect 18924 7586 20668 7588
rect 20764 7586 20870 7702
rect 25990 7696 30348 7704
rect 25990 7688 27316 7696
rect 23282 7686 27316 7688
rect 23282 7684 26922 7686
rect 18924 7582 20870 7586
rect 21270 7680 26922 7684
rect 21270 7678 24996 7680
rect 21270 7670 24524 7678
rect 21270 7668 24104 7670
rect 21270 7658 22682 7668
rect 21270 7646 21748 7658
rect 18924 7580 19452 7582
rect 18234 7576 19452 7580
rect 21270 7574 21406 7646
rect 21506 7574 21748 7646
rect 11276 7570 15412 7574
rect 11276 7564 12772 7570
rect 21270 7564 21748 7574
rect 21884 7654 22682 7658
rect 21884 7582 22242 7654
rect 22342 7582 22682 7654
rect 21884 7574 22682 7582
rect 22818 7666 24104 7668
rect 22818 7594 23152 7666
rect 23252 7594 24104 7666
rect 22818 7580 24104 7594
rect 24216 7588 24524 7670
rect 24636 7590 24996 7678
rect 25108 7670 26922 7680
rect 25108 7590 25442 7670
rect 24636 7588 25442 7590
rect 24216 7580 25442 7588
rect 25554 7668 26922 7670
rect 25554 7580 25886 7668
rect 22818 7578 25886 7580
rect 25998 7584 26922 7668
rect 27028 7594 27316 7686
rect 27422 7690 29436 7696
rect 27422 7676 28278 7690
rect 27422 7594 27776 7676
rect 27028 7584 27776 7594
rect 25998 7578 27776 7584
rect 22818 7576 27776 7578
rect 22818 7574 26020 7576
rect 27882 7588 28278 7676
rect 28384 7676 29436 7690
rect 28384 7588 28736 7676
rect 27882 7576 28736 7588
rect 28842 7580 29436 7676
rect 29532 7682 30348 7696
rect 29532 7590 29856 7682
rect 29946 7590 30348 7682
rect 29532 7588 30348 7590
rect 30444 7702 31478 7704
rect 30444 7684 31276 7702
rect 30444 7592 30802 7684
rect 30892 7592 31276 7684
rect 30444 7588 31276 7592
rect 29532 7586 31276 7588
rect 31372 7586 31478 7702
rect 36518 7696 40876 7704
rect 36518 7688 37844 7696
rect 33810 7686 37844 7688
rect 33810 7684 37450 7686
rect 29532 7582 31478 7586
rect 31798 7680 37450 7684
rect 31798 7678 35524 7680
rect 31798 7670 35052 7678
rect 31798 7668 34632 7670
rect 31798 7658 33210 7668
rect 31798 7646 32276 7658
rect 29532 7580 30060 7582
rect 28842 7576 30060 7580
rect 31798 7574 31934 7646
rect 32034 7574 32276 7646
rect 21884 7570 26020 7574
rect 21884 7564 23380 7570
rect 31798 7564 32276 7574
rect 32412 7654 33210 7658
rect 32412 7582 32770 7654
rect 32870 7582 33210 7654
rect 32412 7574 33210 7582
rect 33346 7666 34632 7668
rect 33346 7594 33680 7666
rect 33780 7594 34632 7666
rect 33346 7580 34632 7594
rect 34744 7588 35052 7670
rect 35164 7590 35524 7678
rect 35636 7670 37450 7680
rect 35636 7590 35970 7670
rect 35164 7588 35970 7590
rect 34744 7580 35970 7588
rect 36082 7668 37450 7670
rect 36082 7580 36414 7668
rect 33346 7578 36414 7580
rect 36526 7584 37450 7668
rect 37556 7594 37844 7686
rect 37950 7690 39964 7696
rect 37950 7676 38806 7690
rect 37950 7594 38304 7676
rect 37556 7584 38304 7594
rect 36526 7578 38304 7584
rect 33346 7576 38304 7578
rect 33346 7574 36548 7576
rect 38410 7588 38806 7676
rect 38912 7676 39964 7690
rect 38912 7588 39264 7676
rect 38410 7576 39264 7588
rect 39370 7580 39964 7676
rect 40060 7682 40876 7696
rect 40060 7590 40384 7682
rect 40474 7590 40876 7682
rect 40060 7588 40876 7590
rect 40972 7702 42006 7704
rect 40972 7684 41804 7702
rect 40972 7592 41330 7684
rect 41420 7592 41804 7684
rect 40972 7588 41804 7592
rect 40060 7586 41804 7588
rect 41900 7586 42006 7702
rect 47128 7696 51486 7704
rect 47128 7688 48454 7696
rect 44420 7686 48454 7688
rect 44420 7684 48060 7686
rect 40060 7582 42006 7586
rect 42408 7680 48060 7684
rect 42408 7678 46134 7680
rect 42408 7670 45662 7678
rect 42408 7668 45242 7670
rect 42408 7658 43820 7668
rect 42408 7646 42886 7658
rect 40060 7580 40588 7582
rect 39370 7576 40588 7580
rect 42408 7574 42544 7646
rect 42644 7574 42886 7646
rect 32412 7570 36548 7574
rect 32412 7564 33908 7570
rect 42408 7564 42886 7574
rect 43022 7654 43820 7658
rect 43022 7582 43380 7654
rect 43480 7582 43820 7654
rect 43022 7574 43820 7582
rect 43956 7666 45242 7668
rect 43956 7594 44290 7666
rect 44390 7594 45242 7666
rect 43956 7580 45242 7594
rect 45354 7588 45662 7670
rect 45774 7590 46134 7678
rect 46246 7670 48060 7680
rect 46246 7590 46580 7670
rect 45774 7588 46580 7590
rect 45354 7580 46580 7588
rect 46692 7668 48060 7670
rect 46692 7580 47024 7668
rect 43956 7578 47024 7580
rect 47136 7584 48060 7668
rect 48166 7594 48454 7686
rect 48560 7690 50574 7696
rect 48560 7676 49416 7690
rect 48560 7594 48914 7676
rect 48166 7584 48914 7594
rect 47136 7578 48914 7584
rect 43956 7576 48914 7578
rect 43956 7574 47158 7576
rect 49020 7588 49416 7676
rect 49522 7676 50574 7690
rect 49522 7588 49874 7676
rect 49020 7576 49874 7588
rect 49980 7580 50574 7676
rect 50670 7682 51486 7696
rect 50670 7590 50994 7682
rect 51084 7590 51486 7682
rect 50670 7588 51486 7590
rect 51582 7702 52616 7704
rect 51582 7684 52414 7702
rect 51582 7592 51940 7684
rect 52030 7592 52414 7684
rect 51582 7588 52414 7592
rect 50670 7586 52414 7588
rect 52510 7586 52616 7702
rect 57656 7696 62014 7704
rect 57656 7688 58982 7696
rect 54948 7686 58982 7688
rect 54948 7684 58588 7686
rect 50670 7582 52616 7586
rect 52936 7680 58588 7684
rect 52936 7678 56662 7680
rect 52936 7670 56190 7678
rect 52936 7668 55770 7670
rect 52936 7658 54348 7668
rect 52936 7646 53414 7658
rect 50670 7580 51198 7582
rect 49980 7576 51198 7580
rect 52936 7574 53072 7646
rect 53172 7574 53414 7646
rect 43022 7570 47158 7574
rect 43022 7564 44518 7570
rect 52936 7564 53414 7574
rect 53550 7654 54348 7658
rect 53550 7582 53908 7654
rect 54008 7582 54348 7654
rect 53550 7574 54348 7582
rect 54484 7666 55770 7668
rect 54484 7594 54818 7666
rect 54918 7594 55770 7666
rect 54484 7580 55770 7594
rect 55882 7588 56190 7670
rect 56302 7590 56662 7678
rect 56774 7670 58588 7680
rect 56774 7590 57108 7670
rect 56302 7588 57108 7590
rect 55882 7580 57108 7588
rect 57220 7668 58588 7670
rect 57220 7580 57552 7668
rect 54484 7578 57552 7580
rect 57664 7584 58588 7668
rect 58694 7594 58982 7686
rect 59088 7690 61102 7696
rect 59088 7676 59944 7690
rect 59088 7594 59442 7676
rect 58694 7584 59442 7594
rect 57664 7578 59442 7584
rect 54484 7576 59442 7578
rect 54484 7574 57686 7576
rect 59548 7588 59944 7676
rect 60050 7676 61102 7690
rect 60050 7588 60402 7676
rect 59548 7576 60402 7588
rect 60508 7580 61102 7676
rect 61198 7682 62014 7696
rect 61198 7590 61522 7682
rect 61612 7590 62014 7682
rect 61198 7588 62014 7590
rect 62110 7702 63144 7704
rect 62110 7684 62942 7702
rect 62110 7592 62468 7684
rect 62558 7592 62942 7684
rect 62110 7588 62942 7592
rect 61198 7586 62942 7588
rect 63038 7586 63144 7702
rect 61198 7582 63144 7586
rect 61198 7580 61726 7582
rect 60508 7576 61726 7580
rect 53550 7570 57686 7574
rect 53550 7564 55046 7570
rect 10646 7386 10742 7394
rect 10646 7360 10732 7386
rect 12644 7360 12740 7394
rect 10646 7298 10680 7360
rect 12706 7298 12740 7360
rect 10806 7258 10822 7292
rect 11190 7258 11206 7292
rect 11264 7258 11280 7292
rect 11648 7258 11664 7292
rect 11722 7258 11738 7292
rect 12106 7258 12122 7292
rect 12180 7258 12196 7292
rect 12564 7258 12580 7292
rect 10760 7199 10794 7215
rect 11218 7199 11252 7215
rect 11676 7199 11710 7215
rect 10760 5207 10794 5223
rect 11218 5207 11252 5223
rect 12134 7199 12168 7215
rect 12592 7199 12626 7215
rect 11676 5207 11710 5223
rect 12134 5207 12168 5223
rect 12592 5207 12626 5223
rect 10806 5161 10822 5164
rect 10806 5130 10815 5161
rect 11190 5130 11206 5164
rect 11264 5161 11280 5164
rect 11264 5130 11273 5161
rect 11648 5130 11664 5164
rect 11722 5161 11738 5164
rect 11722 5130 11731 5161
rect 12106 5130 12122 5164
rect 12180 5161 12196 5164
rect 12180 5130 12189 5161
rect 12564 5130 12580 5164
rect 10646 5062 10680 5124
rect 12706 5062 12740 5124
rect 10646 5028 10742 5062
rect 12644 5028 12740 5062
rect 13400 7354 13496 7388
rect 15398 7354 15494 7388
rect 21254 7386 21350 7394
rect 13400 7292 13434 7354
rect 15460 7292 15494 7354
rect 13560 7252 13576 7286
rect 13944 7252 13960 7286
rect 14018 7252 14034 7286
rect 14402 7252 14418 7286
rect 14476 7252 14492 7286
rect 14860 7252 14876 7286
rect 14934 7252 14950 7286
rect 15318 7252 15334 7286
rect 13514 7193 13548 7209
rect 13972 7193 14006 7209
rect 14430 7193 14464 7209
rect 13514 5201 13548 5217
rect 13972 5201 14006 5217
rect 14430 5201 14464 5217
rect 14888 7193 14922 7209
rect 15346 7193 15380 7209
rect 14888 5201 14922 5217
rect 15346 5201 15380 5217
rect 13560 5124 13576 5158
rect 13944 5124 13960 5158
rect 14018 5124 14034 5158
rect 14402 5124 14418 5158
rect 14476 5124 14492 5158
rect 14860 5124 14876 5158
rect 14934 5124 14950 5158
rect 15318 5124 15334 5158
rect 13400 5056 13434 5118
rect 15460 5056 15494 5118
rect 13400 5022 13496 5056
rect 15398 5022 15494 5056
rect 16216 7328 16312 7362
rect 18214 7328 18310 7362
rect 16216 7266 16250 7328
rect 18276 7266 18310 7328
rect 16376 7226 16392 7260
rect 16760 7226 16776 7260
rect 16834 7226 16850 7260
rect 17218 7226 17234 7260
rect 17292 7226 17308 7260
rect 17676 7226 17692 7260
rect 17750 7226 17766 7260
rect 18134 7226 18150 7260
rect 16330 7167 16364 7183
rect 16788 7167 16822 7183
rect 16330 5175 16364 5191
rect 17246 7167 17280 7183
rect 17704 7167 17738 7183
rect 16788 5175 16822 5191
rect 17246 5175 17280 5191
rect 18162 7167 18196 7183
rect 17704 5175 17738 5191
rect 18162 5175 18196 5191
rect 16376 5098 16392 5132
rect 16760 5098 16776 5132
rect 16834 5098 16850 5132
rect 17218 5098 17234 5132
rect 17292 5098 17308 5132
rect 17676 5098 17692 5132
rect 17750 5098 17766 5132
rect 18134 5098 18150 5132
rect 16216 5030 16250 5092
rect 18276 5030 18310 5092
rect 16216 4996 16312 5030
rect 18214 4996 18310 5030
rect 18740 7350 18836 7384
rect 20738 7350 20834 7384
rect 18740 7288 18774 7350
rect 20800 7288 20834 7350
rect 18900 7248 18916 7282
rect 19284 7248 19300 7282
rect 19358 7248 19374 7282
rect 19742 7248 19758 7282
rect 19816 7248 19832 7282
rect 20200 7248 20216 7282
rect 20274 7248 20290 7282
rect 20658 7248 20674 7282
rect 18854 7189 18888 7205
rect 19312 7189 19346 7205
rect 19770 7189 19804 7205
rect 20228 7189 20262 7205
rect 18854 5197 18888 5213
rect 19312 5197 19346 5213
rect 20686 7189 20720 7205
rect 19770 5197 19804 5213
rect 20228 5197 20262 5213
rect 20686 5197 20720 5213
rect 18900 5120 18916 5154
rect 19284 5120 19300 5154
rect 19358 5120 19374 5154
rect 19742 5120 19758 5154
rect 19816 5120 19832 5154
rect 20200 5120 20216 5154
rect 20274 5120 20290 5154
rect 20658 5120 20674 5154
rect 18740 5052 18774 5114
rect 20800 5052 20834 5114
rect 18740 5018 18836 5052
rect 20738 5018 20834 5052
rect 21254 7360 21340 7386
rect 23252 7360 23348 7394
rect 21254 7298 21288 7360
rect 23314 7298 23348 7360
rect 21414 7258 21430 7292
rect 21798 7258 21814 7292
rect 21872 7258 21888 7292
rect 22256 7258 22272 7292
rect 22330 7258 22346 7292
rect 22714 7258 22730 7292
rect 22788 7258 22804 7292
rect 23172 7258 23188 7292
rect 21368 7199 21402 7215
rect 21826 7199 21860 7215
rect 22284 7199 22318 7215
rect 21368 5207 21402 5223
rect 21826 5207 21860 5223
rect 22742 7199 22776 7215
rect 23200 7199 23234 7215
rect 22284 5207 22318 5223
rect 22742 5207 22776 5223
rect 23200 5207 23234 5223
rect 21414 5161 21430 5164
rect 21414 5130 21423 5161
rect 21798 5130 21814 5164
rect 21872 5161 21888 5164
rect 21872 5130 21881 5161
rect 22256 5130 22272 5164
rect 22330 5161 22346 5164
rect 22330 5130 22339 5161
rect 22714 5130 22730 5164
rect 22788 5161 22804 5164
rect 22788 5130 22797 5161
rect 23172 5130 23188 5164
rect 21254 5062 21288 5124
rect 23314 5062 23348 5124
rect 21254 5028 21350 5062
rect 23252 5028 23348 5062
rect 24008 7354 24104 7388
rect 26006 7354 26102 7388
rect 31782 7386 31878 7394
rect 24008 7292 24042 7354
rect 26068 7292 26102 7354
rect 24168 7252 24184 7286
rect 24552 7252 24568 7286
rect 24626 7252 24642 7286
rect 25010 7252 25026 7286
rect 25084 7252 25100 7286
rect 25468 7252 25484 7286
rect 25542 7252 25558 7286
rect 25926 7252 25942 7286
rect 24122 7193 24156 7209
rect 24580 7193 24614 7209
rect 25038 7193 25072 7209
rect 24122 5201 24156 5217
rect 24580 5201 24614 5217
rect 25038 5201 25072 5217
rect 25496 7193 25530 7209
rect 25954 7193 25988 7209
rect 25496 5201 25530 5217
rect 25954 5201 25988 5217
rect 24168 5124 24184 5158
rect 24552 5124 24568 5158
rect 24626 5124 24642 5158
rect 25010 5124 25026 5158
rect 25084 5124 25100 5158
rect 25468 5124 25484 5158
rect 25542 5124 25558 5158
rect 25926 5124 25942 5158
rect 24008 5056 24042 5118
rect 26068 5056 26102 5118
rect 24008 5022 24104 5056
rect 26006 5022 26102 5056
rect 26824 7328 26920 7362
rect 28822 7328 28918 7362
rect 26824 7266 26858 7328
rect 28884 7266 28918 7328
rect 26984 7226 27000 7260
rect 27368 7226 27384 7260
rect 27442 7226 27458 7260
rect 27826 7226 27842 7260
rect 27900 7226 27916 7260
rect 28284 7226 28300 7260
rect 28358 7226 28374 7260
rect 28742 7226 28758 7260
rect 26938 7167 26972 7183
rect 27396 7167 27430 7183
rect 26938 5175 26972 5191
rect 27854 7167 27888 7183
rect 28312 7167 28346 7183
rect 27396 5175 27430 5191
rect 27854 5175 27888 5191
rect 28770 7167 28804 7183
rect 28312 5175 28346 5191
rect 28770 5175 28804 5191
rect 26984 5098 27000 5132
rect 27368 5098 27384 5132
rect 27442 5098 27458 5132
rect 27826 5098 27842 5132
rect 27900 5098 27916 5132
rect 28284 5098 28300 5132
rect 28358 5098 28374 5132
rect 28742 5098 28758 5132
rect 26824 5030 26858 5092
rect 28884 5030 28918 5092
rect 26824 4996 26920 5030
rect 28822 4996 28918 5030
rect 29348 7350 29444 7384
rect 31346 7350 31442 7384
rect 29348 7288 29382 7350
rect 31408 7288 31442 7350
rect 29508 7248 29524 7282
rect 29892 7248 29908 7282
rect 29966 7248 29982 7282
rect 30350 7248 30366 7282
rect 30424 7248 30440 7282
rect 30808 7248 30824 7282
rect 30882 7248 30898 7282
rect 31266 7248 31282 7282
rect 29462 7189 29496 7205
rect 29920 7189 29954 7205
rect 30378 7189 30412 7205
rect 30836 7189 30870 7205
rect 29462 5197 29496 5213
rect 29920 5197 29954 5213
rect 31294 7189 31328 7205
rect 30378 5197 30412 5213
rect 30836 5197 30870 5213
rect 31294 5197 31328 5213
rect 29508 5120 29524 5154
rect 29892 5120 29908 5154
rect 29966 5120 29982 5154
rect 30350 5120 30366 5154
rect 30424 5120 30440 5154
rect 30808 5120 30824 5154
rect 30882 5120 30898 5154
rect 31266 5120 31282 5154
rect 29348 5052 29382 5114
rect 31408 5052 31442 5114
rect 29348 5018 29444 5052
rect 31346 5018 31442 5052
rect 31782 7360 31868 7386
rect 33780 7360 33876 7394
rect 31782 7298 31816 7360
rect 33842 7298 33876 7360
rect 31942 7258 31958 7292
rect 32326 7258 32342 7292
rect 32400 7258 32416 7292
rect 32784 7258 32800 7292
rect 32858 7258 32874 7292
rect 33242 7258 33258 7292
rect 33316 7258 33332 7292
rect 33700 7258 33716 7292
rect 31896 7199 31930 7215
rect 32354 7199 32388 7215
rect 32812 7199 32846 7215
rect 31896 5207 31930 5223
rect 32354 5207 32388 5223
rect 33270 7199 33304 7215
rect 33728 7199 33762 7215
rect 32812 5207 32846 5223
rect 33270 5207 33304 5223
rect 33728 5207 33762 5223
rect 31942 5161 31958 5164
rect 31942 5130 31951 5161
rect 32326 5130 32342 5164
rect 32400 5161 32416 5164
rect 32400 5130 32409 5161
rect 32784 5130 32800 5164
rect 32858 5161 32874 5164
rect 32858 5130 32867 5161
rect 33242 5130 33258 5164
rect 33316 5161 33332 5164
rect 33316 5130 33325 5161
rect 33700 5130 33716 5164
rect 31782 5062 31816 5124
rect 33842 5062 33876 5124
rect 31782 5028 31878 5062
rect 33780 5028 33876 5062
rect 34536 7354 34632 7388
rect 36534 7354 36630 7388
rect 42392 7386 42488 7394
rect 34536 7292 34570 7354
rect 36596 7292 36630 7354
rect 34696 7252 34712 7286
rect 35080 7252 35096 7286
rect 35154 7252 35170 7286
rect 35538 7252 35554 7286
rect 35612 7252 35628 7286
rect 35996 7252 36012 7286
rect 36070 7252 36086 7286
rect 36454 7252 36470 7286
rect 34650 7193 34684 7209
rect 35108 7193 35142 7209
rect 35566 7193 35600 7209
rect 34650 5201 34684 5217
rect 35108 5201 35142 5217
rect 35566 5201 35600 5217
rect 36024 7193 36058 7209
rect 36482 7193 36516 7209
rect 36024 5201 36058 5217
rect 36482 5201 36516 5217
rect 34696 5124 34712 5158
rect 35080 5124 35096 5158
rect 35154 5124 35170 5158
rect 35538 5124 35554 5158
rect 35612 5124 35628 5158
rect 35996 5124 36012 5158
rect 36070 5124 36086 5158
rect 36454 5124 36470 5158
rect 34536 5056 34570 5118
rect 36596 5056 36630 5118
rect 34536 5022 34632 5056
rect 36534 5022 36630 5056
rect 37352 7328 37448 7362
rect 39350 7328 39446 7362
rect 37352 7266 37386 7328
rect 39412 7266 39446 7328
rect 37512 7226 37528 7260
rect 37896 7226 37912 7260
rect 37970 7226 37986 7260
rect 38354 7226 38370 7260
rect 38428 7226 38444 7260
rect 38812 7226 38828 7260
rect 38886 7226 38902 7260
rect 39270 7226 39286 7260
rect 37466 7167 37500 7183
rect 37924 7167 37958 7183
rect 37466 5175 37500 5191
rect 38382 7167 38416 7183
rect 38840 7167 38874 7183
rect 37924 5175 37958 5191
rect 38382 5175 38416 5191
rect 39298 7167 39332 7183
rect 38840 5175 38874 5191
rect 39298 5175 39332 5191
rect 37512 5098 37528 5132
rect 37896 5098 37912 5132
rect 37970 5098 37986 5132
rect 38354 5098 38370 5132
rect 38428 5098 38444 5132
rect 38812 5098 38828 5132
rect 38886 5098 38902 5132
rect 39270 5098 39286 5132
rect 37352 5030 37386 5092
rect 39412 5030 39446 5092
rect 37352 4996 37448 5030
rect 39350 4996 39446 5030
rect 39876 7350 39972 7384
rect 41874 7350 41970 7384
rect 39876 7288 39910 7350
rect 41936 7288 41970 7350
rect 40036 7248 40052 7282
rect 40420 7248 40436 7282
rect 40494 7248 40510 7282
rect 40878 7248 40894 7282
rect 40952 7248 40968 7282
rect 41336 7248 41352 7282
rect 41410 7248 41426 7282
rect 41794 7248 41810 7282
rect 39990 7189 40024 7205
rect 40448 7189 40482 7205
rect 40906 7189 40940 7205
rect 41364 7189 41398 7205
rect 39990 5197 40024 5213
rect 40448 5197 40482 5213
rect 41822 7189 41856 7205
rect 40906 5197 40940 5213
rect 41364 5197 41398 5213
rect 41822 5197 41856 5213
rect 40036 5120 40052 5154
rect 40420 5120 40436 5154
rect 40494 5120 40510 5154
rect 40878 5120 40894 5154
rect 40952 5120 40968 5154
rect 41336 5120 41352 5154
rect 41410 5120 41426 5154
rect 41794 5120 41810 5154
rect 39876 5052 39910 5114
rect 41936 5052 41970 5114
rect 39876 5018 39972 5052
rect 41874 5018 41970 5052
rect 42392 7360 42478 7386
rect 44390 7360 44486 7394
rect 42392 7298 42426 7360
rect 44452 7298 44486 7360
rect 42552 7258 42568 7292
rect 42936 7258 42952 7292
rect 43010 7258 43026 7292
rect 43394 7258 43410 7292
rect 43468 7258 43484 7292
rect 43852 7258 43868 7292
rect 43926 7258 43942 7292
rect 44310 7258 44326 7292
rect 42506 7199 42540 7215
rect 42964 7199 42998 7215
rect 43422 7199 43456 7215
rect 42506 5207 42540 5223
rect 42964 5207 42998 5223
rect 43880 7199 43914 7215
rect 44338 7199 44372 7215
rect 43422 5207 43456 5223
rect 43880 5207 43914 5223
rect 44338 5207 44372 5223
rect 42552 5161 42568 5164
rect 42552 5130 42561 5161
rect 42936 5130 42952 5164
rect 43010 5161 43026 5164
rect 43010 5130 43019 5161
rect 43394 5130 43410 5164
rect 43468 5161 43484 5164
rect 43468 5130 43477 5161
rect 43852 5130 43868 5164
rect 43926 5161 43942 5164
rect 43926 5130 43935 5161
rect 44310 5130 44326 5164
rect 42392 5062 42426 5124
rect 44452 5062 44486 5124
rect 42392 5028 42488 5062
rect 44390 5028 44486 5062
rect 45146 7354 45242 7388
rect 47144 7354 47240 7388
rect 52920 7386 53016 7394
rect 45146 7292 45180 7354
rect 47206 7292 47240 7354
rect 45306 7252 45322 7286
rect 45690 7252 45706 7286
rect 45764 7252 45780 7286
rect 46148 7252 46164 7286
rect 46222 7252 46238 7286
rect 46606 7252 46622 7286
rect 46680 7252 46696 7286
rect 47064 7252 47080 7286
rect 45260 7193 45294 7209
rect 45718 7193 45752 7209
rect 46176 7193 46210 7209
rect 45260 5201 45294 5217
rect 45718 5201 45752 5217
rect 46176 5201 46210 5217
rect 46634 7193 46668 7209
rect 47092 7193 47126 7209
rect 46634 5201 46668 5217
rect 47092 5201 47126 5217
rect 45306 5124 45322 5158
rect 45690 5124 45706 5158
rect 45764 5124 45780 5158
rect 46148 5124 46164 5158
rect 46222 5124 46238 5158
rect 46606 5124 46622 5158
rect 46680 5124 46696 5158
rect 47064 5124 47080 5158
rect 45146 5056 45180 5118
rect 47206 5056 47240 5118
rect 45146 5022 45242 5056
rect 47144 5022 47240 5056
rect 47962 7328 48058 7362
rect 49960 7328 50056 7362
rect 47962 7266 47996 7328
rect 50022 7266 50056 7328
rect 48122 7226 48138 7260
rect 48506 7226 48522 7260
rect 48580 7226 48596 7260
rect 48964 7226 48980 7260
rect 49038 7226 49054 7260
rect 49422 7226 49438 7260
rect 49496 7226 49512 7260
rect 49880 7226 49896 7260
rect 48076 7167 48110 7183
rect 48534 7167 48568 7183
rect 48076 5175 48110 5191
rect 48992 7167 49026 7183
rect 49450 7167 49484 7183
rect 48534 5175 48568 5191
rect 48992 5175 49026 5191
rect 49908 7167 49942 7183
rect 49450 5175 49484 5191
rect 49908 5175 49942 5191
rect 48122 5098 48138 5132
rect 48506 5098 48522 5132
rect 48580 5098 48596 5132
rect 48964 5098 48980 5132
rect 49038 5098 49054 5132
rect 49422 5098 49438 5132
rect 49496 5098 49512 5132
rect 49880 5098 49896 5132
rect 47962 5030 47996 5092
rect 50022 5030 50056 5092
rect 47962 4996 48058 5030
rect 49960 4996 50056 5030
rect 50486 7350 50582 7384
rect 52484 7350 52580 7384
rect 50486 7288 50520 7350
rect 52546 7288 52580 7350
rect 50646 7248 50662 7282
rect 51030 7248 51046 7282
rect 51104 7248 51120 7282
rect 51488 7248 51504 7282
rect 51562 7248 51578 7282
rect 51946 7248 51962 7282
rect 52020 7248 52036 7282
rect 52404 7248 52420 7282
rect 50600 7189 50634 7205
rect 51058 7189 51092 7205
rect 51516 7189 51550 7205
rect 51974 7189 52008 7205
rect 50600 5197 50634 5213
rect 51058 5197 51092 5213
rect 52432 7189 52466 7205
rect 51516 5197 51550 5213
rect 51974 5197 52008 5213
rect 52432 5197 52466 5213
rect 50646 5120 50662 5154
rect 51030 5120 51046 5154
rect 51104 5120 51120 5154
rect 51488 5120 51504 5154
rect 51562 5120 51578 5154
rect 51946 5120 51962 5154
rect 52020 5120 52036 5154
rect 52404 5120 52420 5154
rect 50486 5052 50520 5114
rect 52546 5052 52580 5114
rect 50486 5018 50582 5052
rect 52484 5018 52580 5052
rect 52920 7360 53006 7386
rect 54918 7360 55014 7394
rect 52920 7298 52954 7360
rect 54980 7298 55014 7360
rect 53080 7258 53096 7292
rect 53464 7258 53480 7292
rect 53538 7258 53554 7292
rect 53922 7258 53938 7292
rect 53996 7258 54012 7292
rect 54380 7258 54396 7292
rect 54454 7258 54470 7292
rect 54838 7258 54854 7292
rect 53034 7199 53068 7215
rect 53492 7199 53526 7215
rect 53950 7199 53984 7215
rect 53034 5207 53068 5223
rect 53492 5207 53526 5223
rect 54408 7199 54442 7215
rect 54866 7199 54900 7215
rect 53950 5207 53984 5223
rect 54408 5207 54442 5223
rect 54866 5207 54900 5223
rect 53080 5161 53096 5164
rect 53080 5130 53089 5161
rect 53464 5130 53480 5164
rect 53538 5161 53554 5164
rect 53538 5130 53547 5161
rect 53922 5130 53938 5164
rect 53996 5161 54012 5164
rect 53996 5130 54005 5161
rect 54380 5130 54396 5164
rect 54454 5161 54470 5164
rect 54454 5130 54463 5161
rect 54838 5130 54854 5164
rect 52920 5062 52954 5124
rect 54980 5062 55014 5124
rect 52920 5028 53016 5062
rect 54918 5028 55014 5062
rect 55674 7354 55770 7388
rect 57672 7354 57768 7388
rect 55674 7292 55708 7354
rect 57734 7292 57768 7354
rect 55834 7252 55850 7286
rect 56218 7252 56234 7286
rect 56292 7252 56308 7286
rect 56676 7252 56692 7286
rect 56750 7252 56766 7286
rect 57134 7252 57150 7286
rect 57208 7252 57224 7286
rect 57592 7252 57608 7286
rect 55788 7193 55822 7209
rect 56246 7193 56280 7209
rect 56704 7193 56738 7209
rect 55788 5201 55822 5217
rect 56246 5201 56280 5217
rect 56704 5201 56738 5217
rect 57162 7193 57196 7209
rect 57620 7193 57654 7209
rect 57162 5201 57196 5217
rect 57620 5201 57654 5217
rect 55834 5124 55850 5158
rect 56218 5124 56234 5158
rect 56292 5124 56308 5158
rect 56676 5124 56692 5158
rect 56750 5124 56766 5158
rect 57134 5124 57150 5158
rect 57208 5124 57224 5158
rect 57592 5124 57608 5158
rect 55674 5056 55708 5118
rect 57734 5056 57768 5118
rect 55674 5022 55770 5056
rect 57672 5022 57768 5056
rect 58490 7328 58586 7362
rect 60488 7328 60584 7362
rect 58490 7266 58524 7328
rect 60550 7266 60584 7328
rect 58650 7226 58666 7260
rect 59034 7226 59050 7260
rect 59108 7226 59124 7260
rect 59492 7226 59508 7260
rect 59566 7226 59582 7260
rect 59950 7226 59966 7260
rect 60024 7226 60040 7260
rect 60408 7226 60424 7260
rect 58604 7167 58638 7183
rect 59062 7167 59096 7183
rect 58604 5175 58638 5191
rect 59520 7167 59554 7183
rect 59978 7167 60012 7183
rect 59062 5175 59096 5191
rect 59520 5175 59554 5191
rect 60436 7167 60470 7183
rect 59978 5175 60012 5191
rect 60436 5175 60470 5191
rect 58650 5098 58666 5132
rect 59034 5098 59050 5132
rect 59108 5098 59124 5132
rect 59492 5098 59508 5132
rect 59566 5098 59582 5132
rect 59950 5098 59966 5132
rect 60024 5098 60040 5132
rect 60408 5098 60424 5132
rect 58490 5030 58524 5092
rect 60550 5030 60584 5092
rect 58490 4996 58586 5030
rect 60488 4996 60584 5030
rect 61014 7350 61110 7384
rect 63012 7350 63108 7384
rect 61014 7288 61048 7350
rect 63074 7288 63108 7350
rect 61174 7248 61190 7282
rect 61558 7248 61574 7282
rect 61632 7248 61648 7282
rect 62016 7248 62032 7282
rect 62090 7248 62106 7282
rect 62474 7248 62490 7282
rect 62548 7248 62564 7282
rect 62932 7248 62948 7282
rect 61128 7189 61162 7205
rect 61586 7189 61620 7205
rect 62044 7189 62078 7205
rect 62502 7189 62536 7205
rect 61128 5197 61162 5213
rect 61586 5197 61620 5213
rect 62960 7189 62994 7205
rect 62044 5197 62078 5213
rect 62502 5197 62536 5213
rect 62960 5197 62994 5213
rect 61174 5120 61190 5154
rect 61558 5120 61574 5154
rect 61632 5120 61648 5154
rect 62016 5120 62032 5154
rect 62090 5120 62106 5154
rect 62474 5120 62490 5154
rect 62548 5120 62564 5154
rect 62932 5120 62948 5154
rect 61014 5052 61048 5114
rect 63074 5052 63108 5114
rect 61014 5018 61110 5052
rect 63012 5018 63108 5052
rect 11906 4202 12002 4236
rect 14158 4202 14254 4236
rect 11906 4140 11940 4202
rect 14220 4140 14254 4202
rect 12008 4078 12042 4094
rect 12076 4088 12092 4122
rect 14068 4088 14084 4122
rect 12008 4028 12042 4044
rect 14118 4078 14152 4094
rect 12076 4000 12092 4034
rect 14068 4000 14084 4034
rect 14118 4028 14152 4044
rect 11906 3920 11940 3982
rect 14220 3920 14254 3982
rect 11906 3886 12002 3920
rect 14158 3886 14254 3920
rect 17356 4212 17452 4246
rect 19608 4212 19704 4246
rect 17356 4150 17390 4212
rect 19670 4150 19704 4212
rect 17458 4088 17492 4104
rect 17526 4098 17542 4132
rect 19518 4098 19534 4132
rect 17458 4038 17492 4054
rect 19568 4088 19602 4104
rect 17526 4010 17542 4044
rect 19518 4010 19534 4044
rect 19568 4038 19602 4054
rect 17356 3930 17390 3992
rect 19670 3930 19704 3992
rect 17356 3896 17452 3930
rect 19608 3896 19704 3930
rect 22514 4202 22610 4236
rect 24766 4202 24862 4236
rect 22514 4140 22548 4202
rect 24828 4140 24862 4202
rect 22616 4078 22650 4094
rect 22684 4088 22700 4122
rect 24676 4088 24692 4122
rect 22616 4028 22650 4044
rect 24726 4078 24760 4094
rect 22684 4000 22700 4034
rect 24676 4000 24692 4034
rect 24726 4028 24760 4044
rect 22514 3920 22548 3982
rect 24828 3920 24862 3982
rect 22514 3886 22610 3920
rect 24766 3886 24862 3920
rect 27964 4212 28060 4246
rect 30216 4212 30312 4246
rect 27964 4150 27998 4212
rect 30278 4150 30312 4212
rect 28066 4088 28100 4104
rect 28134 4098 28150 4132
rect 30126 4098 30142 4132
rect 28066 4038 28100 4054
rect 30176 4088 30210 4104
rect 28134 4010 28150 4044
rect 30126 4010 30142 4044
rect 30176 4038 30210 4054
rect 27964 3930 27998 3992
rect 30278 3930 30312 3992
rect 27964 3896 28060 3930
rect 30216 3896 30312 3930
rect 33042 4202 33138 4236
rect 35294 4202 35390 4236
rect 33042 4140 33076 4202
rect 35356 4140 35390 4202
rect 33144 4078 33178 4094
rect 33212 4088 33228 4122
rect 35204 4088 35220 4122
rect 33144 4028 33178 4044
rect 35254 4078 35288 4094
rect 33212 4000 33228 4034
rect 35204 4000 35220 4034
rect 35254 4028 35288 4044
rect 33042 3920 33076 3982
rect 35356 3920 35390 3982
rect 33042 3886 33138 3920
rect 35294 3886 35390 3920
rect 38492 4212 38588 4246
rect 40744 4212 40840 4246
rect 38492 4150 38526 4212
rect 40806 4150 40840 4212
rect 38594 4088 38628 4104
rect 38662 4098 38678 4132
rect 40654 4098 40670 4132
rect 38594 4038 38628 4054
rect 40704 4088 40738 4104
rect 38662 4010 38678 4044
rect 40654 4010 40670 4044
rect 40704 4038 40738 4054
rect 38492 3930 38526 3992
rect 40806 3930 40840 3992
rect 38492 3896 38588 3930
rect 40744 3896 40840 3930
rect 43652 4202 43748 4236
rect 45904 4202 46000 4236
rect 43652 4140 43686 4202
rect 45966 4140 46000 4202
rect 43754 4078 43788 4094
rect 43822 4088 43838 4122
rect 45814 4088 45830 4122
rect 43754 4028 43788 4044
rect 45864 4078 45898 4094
rect 43822 4000 43838 4034
rect 45814 4000 45830 4034
rect 45864 4028 45898 4044
rect 43652 3920 43686 3982
rect 45966 3920 46000 3982
rect 43652 3886 43748 3920
rect 45904 3886 46000 3920
rect 49102 4212 49198 4246
rect 51354 4212 51450 4246
rect 49102 4150 49136 4212
rect 51416 4150 51450 4212
rect 49204 4088 49238 4104
rect 49272 4098 49288 4132
rect 51264 4098 51280 4132
rect 49204 4038 49238 4054
rect 51314 4088 51348 4104
rect 49272 4010 49288 4044
rect 51264 4010 51280 4044
rect 51314 4038 51348 4054
rect 49102 3930 49136 3992
rect 51416 3930 51450 3992
rect 49102 3896 49198 3930
rect 51354 3896 51450 3930
rect 54180 4202 54276 4236
rect 56432 4202 56528 4236
rect 54180 4140 54214 4202
rect 56494 4140 56528 4202
rect 54282 4078 54316 4094
rect 54350 4088 54366 4122
rect 56342 4088 56358 4122
rect 54282 4028 54316 4044
rect 56392 4078 56426 4094
rect 54350 4000 54366 4034
rect 56342 4000 56358 4034
rect 56392 4028 56426 4044
rect 54180 3920 54214 3982
rect 56494 3920 56528 3982
rect 54180 3886 54276 3920
rect 56432 3886 56528 3920
rect 59630 4212 59726 4246
rect 61882 4212 61978 4246
rect 59630 4150 59664 4212
rect 61944 4150 61978 4212
rect 59732 4088 59766 4104
rect 59800 4098 59816 4132
rect 61792 4098 61808 4132
rect 59732 4038 59766 4054
rect 61842 4088 61876 4104
rect 59800 4010 59816 4044
rect 61792 4010 61808 4044
rect 61842 4038 61876 4054
rect 59630 3930 59664 3992
rect 61944 3930 61978 3992
rect 59630 3896 59726 3930
rect 61882 3896 61978 3930
rect 14315 3193 14411 3227
rect 19519 3193 19615 3227
rect 14315 3131 14349 3193
rect 19581 3131 19615 3193
rect 14475 3091 14491 3125
rect 14859 3091 14875 3125
rect 14933 3091 14949 3125
rect 15317 3091 15333 3125
rect 15391 3091 15407 3125
rect 15775 3091 15791 3125
rect 15849 3091 15865 3125
rect 16233 3091 16249 3125
rect 16307 3091 16323 3125
rect 16691 3091 16707 3125
rect 16765 3091 16781 3125
rect 17149 3091 17165 3125
rect 17223 3091 17239 3125
rect 17607 3091 17623 3125
rect 17681 3091 17697 3125
rect 18065 3091 18081 3125
rect 18139 3091 18155 3125
rect 18523 3091 18539 3125
rect 18597 3091 18613 3125
rect 18981 3091 18997 3125
rect 19055 3091 19071 3125
rect 19439 3091 19455 3125
rect 14429 3041 14463 3057
rect 14887 3041 14921 3057
rect 15345 3041 15379 3057
rect 15803 3041 15837 3057
rect 14429 649 14463 665
rect 14887 649 14921 665
rect 16261 3041 16295 3057
rect 16719 3041 16753 3057
rect 15345 649 15379 665
rect 15803 649 15837 665
rect 17177 3041 17211 3057
rect 17635 3041 17669 3057
rect 16261 649 16295 665
rect 16719 649 16753 665
rect 18093 3041 18127 3057
rect 17177 649 17211 665
rect 17635 649 17669 665
rect 18551 3041 18585 3057
rect 19009 3041 19043 3057
rect 19467 3041 19501 3057
rect 18093 649 18127 665
rect 18551 649 18585 665
rect 19009 649 19043 665
rect 19467 649 19501 665
rect 14475 581 14491 615
rect 14859 581 14875 615
rect 14933 581 14949 615
rect 15317 581 15333 615
rect 15391 581 15407 615
rect 15775 581 15791 615
rect 15849 581 15865 615
rect 16233 581 16249 615
rect 16307 581 16323 615
rect 16691 581 16707 615
rect 16765 581 16781 615
rect 17149 581 17165 615
rect 17223 581 17239 615
rect 17607 581 17623 615
rect 17681 581 17697 615
rect 18065 581 18081 615
rect 18139 581 18155 615
rect 18523 581 18539 615
rect 18597 581 18613 615
rect 18981 581 18997 615
rect 19055 581 19071 615
rect 19439 581 19455 615
rect 14315 513 14349 575
rect 19581 513 19615 575
rect 14315 479 14411 513
rect 19519 479 19615 513
rect 24923 3193 25019 3227
rect 30127 3193 30223 3227
rect 24923 3131 24957 3193
rect 30189 3131 30223 3193
rect 25083 3091 25099 3125
rect 25467 3091 25483 3125
rect 25541 3091 25557 3125
rect 25925 3091 25941 3125
rect 25999 3091 26015 3125
rect 26383 3091 26399 3125
rect 26457 3091 26473 3125
rect 26841 3091 26857 3125
rect 26915 3091 26931 3125
rect 27299 3091 27315 3125
rect 27373 3091 27389 3125
rect 27757 3091 27773 3125
rect 27831 3091 27847 3125
rect 28215 3091 28231 3125
rect 28289 3091 28305 3125
rect 28673 3091 28689 3125
rect 28747 3091 28763 3125
rect 29131 3091 29147 3125
rect 29205 3091 29221 3125
rect 29589 3091 29605 3125
rect 29663 3091 29679 3125
rect 30047 3091 30063 3125
rect 25037 3041 25071 3057
rect 25495 3041 25529 3057
rect 25953 3041 25987 3057
rect 26411 3041 26445 3057
rect 25037 649 25071 665
rect 25495 649 25529 665
rect 26869 3041 26903 3057
rect 27327 3041 27361 3057
rect 25953 649 25987 665
rect 26411 649 26445 665
rect 27785 3041 27819 3057
rect 28243 3041 28277 3057
rect 26869 649 26903 665
rect 27327 649 27361 665
rect 28701 3041 28735 3057
rect 27785 649 27819 665
rect 28243 649 28277 665
rect 29159 3041 29193 3057
rect 29617 3041 29651 3057
rect 30075 3041 30109 3057
rect 28701 649 28735 665
rect 29159 649 29193 665
rect 29617 649 29651 665
rect 30075 649 30109 665
rect 25083 581 25099 615
rect 25467 581 25483 615
rect 25541 581 25557 615
rect 25925 581 25941 615
rect 25999 581 26015 615
rect 26383 581 26399 615
rect 26457 581 26473 615
rect 26841 581 26857 615
rect 26915 581 26931 615
rect 27299 581 27315 615
rect 27373 581 27389 615
rect 27757 581 27773 615
rect 27831 581 27847 615
rect 28215 581 28231 615
rect 28289 581 28305 615
rect 28673 581 28689 615
rect 28747 581 28763 615
rect 29131 581 29147 615
rect 29205 581 29221 615
rect 29589 581 29605 615
rect 29663 581 29679 615
rect 30047 581 30063 615
rect 24923 513 24957 575
rect 30189 513 30223 575
rect 24923 479 25019 513
rect 30127 479 30223 513
rect 35451 3193 35547 3227
rect 40655 3193 40751 3227
rect 35451 3131 35485 3193
rect 40717 3131 40751 3193
rect 35611 3091 35627 3125
rect 35995 3091 36011 3125
rect 36069 3091 36085 3125
rect 36453 3091 36469 3125
rect 36527 3091 36543 3125
rect 36911 3091 36927 3125
rect 36985 3091 37001 3125
rect 37369 3091 37385 3125
rect 37443 3091 37459 3125
rect 37827 3091 37843 3125
rect 37901 3091 37917 3125
rect 38285 3091 38301 3125
rect 38359 3091 38375 3125
rect 38743 3091 38759 3125
rect 38817 3091 38833 3125
rect 39201 3091 39217 3125
rect 39275 3091 39291 3125
rect 39659 3091 39675 3125
rect 39733 3091 39749 3125
rect 40117 3091 40133 3125
rect 40191 3091 40207 3125
rect 40575 3091 40591 3125
rect 35565 3041 35599 3057
rect 36023 3041 36057 3057
rect 36481 3041 36515 3057
rect 36939 3041 36973 3057
rect 35565 649 35599 665
rect 36023 649 36057 665
rect 37397 3041 37431 3057
rect 37855 3041 37889 3057
rect 36481 649 36515 665
rect 36939 649 36973 665
rect 38313 3041 38347 3057
rect 38771 3041 38805 3057
rect 37397 649 37431 665
rect 37855 649 37889 665
rect 39229 3041 39263 3057
rect 38313 649 38347 665
rect 38771 649 38805 665
rect 39687 3041 39721 3057
rect 40145 3041 40179 3057
rect 40603 3041 40637 3057
rect 39229 649 39263 665
rect 39687 649 39721 665
rect 40145 649 40179 665
rect 40603 649 40637 665
rect 35611 581 35627 615
rect 35995 581 36011 615
rect 36069 581 36085 615
rect 36453 581 36469 615
rect 36527 581 36543 615
rect 36911 581 36927 615
rect 36985 581 37001 615
rect 37369 581 37385 615
rect 37443 581 37459 615
rect 37827 581 37843 615
rect 37901 581 37917 615
rect 38285 581 38301 615
rect 38359 581 38375 615
rect 38743 581 38759 615
rect 38817 581 38833 615
rect 39201 581 39217 615
rect 39275 581 39291 615
rect 39659 581 39675 615
rect 39733 581 39749 615
rect 40117 581 40133 615
rect 40191 581 40207 615
rect 40575 581 40591 615
rect 35451 513 35485 575
rect 40717 513 40751 575
rect 35451 479 35547 513
rect 40655 479 40751 513
rect 46061 3193 46157 3227
rect 51265 3193 51361 3227
rect 46061 3131 46095 3193
rect 51327 3131 51361 3193
rect 46221 3091 46237 3125
rect 46605 3091 46621 3125
rect 46679 3091 46695 3125
rect 47063 3091 47079 3125
rect 47137 3091 47153 3125
rect 47521 3091 47537 3125
rect 47595 3091 47611 3125
rect 47979 3091 47995 3125
rect 48053 3091 48069 3125
rect 48437 3091 48453 3125
rect 48511 3091 48527 3125
rect 48895 3091 48911 3125
rect 48969 3091 48985 3125
rect 49353 3091 49369 3125
rect 49427 3091 49443 3125
rect 49811 3091 49827 3125
rect 49885 3091 49901 3125
rect 50269 3091 50285 3125
rect 50343 3091 50359 3125
rect 50727 3091 50743 3125
rect 50801 3091 50817 3125
rect 51185 3091 51201 3125
rect 46175 3041 46209 3057
rect 46633 3041 46667 3057
rect 47091 3041 47125 3057
rect 47549 3041 47583 3057
rect 46175 649 46209 665
rect 46633 649 46667 665
rect 48007 3041 48041 3057
rect 48465 3041 48499 3057
rect 47091 649 47125 665
rect 47549 649 47583 665
rect 48923 3041 48957 3057
rect 49381 3041 49415 3057
rect 48007 649 48041 665
rect 48465 649 48499 665
rect 49839 3041 49873 3057
rect 48923 649 48957 665
rect 49381 649 49415 665
rect 50297 3041 50331 3057
rect 50755 3041 50789 3057
rect 51213 3041 51247 3057
rect 49839 649 49873 665
rect 50297 649 50331 665
rect 50755 649 50789 665
rect 51213 649 51247 665
rect 46221 581 46237 615
rect 46605 581 46621 615
rect 46679 581 46695 615
rect 47063 581 47079 615
rect 47137 581 47153 615
rect 47521 581 47537 615
rect 47595 581 47611 615
rect 47979 581 47995 615
rect 48053 581 48069 615
rect 48437 581 48453 615
rect 48511 581 48527 615
rect 48895 581 48911 615
rect 48969 581 48985 615
rect 49353 581 49369 615
rect 49427 581 49443 615
rect 49811 581 49827 615
rect 49885 581 49901 615
rect 50269 581 50285 615
rect 50343 581 50359 615
rect 50727 581 50743 615
rect 50801 581 50817 615
rect 51185 581 51201 615
rect 46061 513 46095 575
rect 51327 513 51361 575
rect 46061 479 46157 513
rect 51265 479 51361 513
rect 56589 3193 56685 3227
rect 61793 3193 61889 3227
rect 56589 3131 56623 3193
rect 61855 3131 61889 3193
rect 56749 3091 56765 3125
rect 57133 3091 57149 3125
rect 57207 3091 57223 3125
rect 57591 3091 57607 3125
rect 57665 3091 57681 3125
rect 58049 3091 58065 3125
rect 58123 3091 58139 3125
rect 58507 3091 58523 3125
rect 58581 3091 58597 3125
rect 58965 3091 58981 3125
rect 59039 3091 59055 3125
rect 59423 3091 59439 3125
rect 59497 3091 59513 3125
rect 59881 3091 59897 3125
rect 59955 3091 59971 3125
rect 60339 3091 60355 3125
rect 60413 3091 60429 3125
rect 60797 3091 60813 3125
rect 60871 3091 60887 3125
rect 61255 3091 61271 3125
rect 61329 3091 61345 3125
rect 61713 3091 61729 3125
rect 56703 3041 56737 3057
rect 57161 3041 57195 3057
rect 57619 3041 57653 3057
rect 58077 3041 58111 3057
rect 56703 649 56737 665
rect 57161 649 57195 665
rect 58535 3041 58569 3057
rect 58993 3041 59027 3057
rect 57619 649 57653 665
rect 58077 649 58111 665
rect 59451 3041 59485 3057
rect 59909 3041 59943 3057
rect 58535 649 58569 665
rect 58993 649 59027 665
rect 60367 3041 60401 3057
rect 59451 649 59485 665
rect 59909 649 59943 665
rect 60825 3041 60859 3057
rect 61283 3041 61317 3057
rect 61741 3041 61775 3057
rect 60367 649 60401 665
rect 60825 649 60859 665
rect 61283 649 61317 665
rect 61741 649 61775 665
rect 56749 581 56765 615
rect 57133 581 57149 615
rect 57207 581 57223 615
rect 57591 581 57607 615
rect 57665 581 57681 615
rect 58049 581 58065 615
rect 58123 581 58139 615
rect 58507 581 58523 615
rect 58581 581 58597 615
rect 58965 581 58981 615
rect 59039 581 59055 615
rect 59423 581 59439 615
rect 59497 581 59513 615
rect 59881 581 59897 615
rect 59955 581 59971 615
rect 60339 581 60355 615
rect 60413 581 60429 615
rect 60797 581 60813 615
rect 60871 581 60887 615
rect 61255 581 61271 615
rect 61329 581 61345 615
rect 61713 581 61729 615
rect 56589 513 56623 575
rect 61855 513 61889 575
rect 56589 479 56685 513
rect 61793 479 61889 513
rect 14270 278 19748 280
rect 14270 272 17148 278
rect 14270 164 14372 272
rect 14486 264 16208 272
rect 14486 258 15722 264
rect 14486 164 14828 258
rect 14270 142 14828 164
rect 14986 256 15722 258
rect 14986 148 15318 256
rect 15432 148 15722 256
rect 15880 164 16208 264
rect 16322 170 17148 272
rect 17262 272 18970 278
rect 17262 264 18076 272
rect 17262 170 17492 264
rect 16322 164 17492 170
rect 15880 148 17492 164
rect 17650 164 18076 264
rect 18190 268 18970 272
rect 18190 164 18590 268
rect 17650 152 18590 164
rect 18748 170 18970 268
rect 19084 170 19748 278
rect 18748 152 19748 170
rect 17650 148 19748 152
rect 14986 142 19748 148
rect 14270 130 19748 142
rect 24878 278 30356 280
rect 24878 272 27756 278
rect 24878 164 24980 272
rect 25094 264 26816 272
rect 25094 258 26330 264
rect 25094 164 25436 258
rect 24878 142 25436 164
rect 25594 256 26330 258
rect 25594 148 25926 256
rect 26040 148 26330 256
rect 26488 164 26816 264
rect 26930 170 27756 272
rect 27870 272 29578 278
rect 27870 264 28684 272
rect 27870 170 28100 264
rect 26930 164 28100 170
rect 26488 148 28100 164
rect 28258 164 28684 264
rect 28798 268 29578 272
rect 28798 164 29198 268
rect 28258 152 29198 164
rect 29356 170 29578 268
rect 29692 170 30356 278
rect 29356 152 30356 170
rect 28258 148 30356 152
rect 25594 142 30356 148
rect 24878 130 30356 142
rect 35406 278 40884 280
rect 35406 272 38284 278
rect 35406 164 35508 272
rect 35622 264 37344 272
rect 35622 258 36858 264
rect 35622 164 35964 258
rect 35406 142 35964 164
rect 36122 256 36858 258
rect 36122 148 36454 256
rect 36568 148 36858 256
rect 37016 164 37344 264
rect 37458 170 38284 272
rect 38398 272 40106 278
rect 38398 264 39212 272
rect 38398 170 38628 264
rect 37458 164 38628 170
rect 37016 148 38628 164
rect 38786 164 39212 264
rect 39326 268 40106 272
rect 39326 164 39726 268
rect 38786 152 39726 164
rect 39884 170 40106 268
rect 40220 170 40884 278
rect 39884 152 40884 170
rect 38786 148 40884 152
rect 36122 142 40884 148
rect 35406 130 40884 142
rect 46016 278 51494 280
rect 46016 272 48894 278
rect 46016 164 46118 272
rect 46232 264 47954 272
rect 46232 258 47468 264
rect 46232 164 46574 258
rect 46016 142 46574 164
rect 46732 256 47468 258
rect 46732 148 47064 256
rect 47178 148 47468 256
rect 47626 164 47954 264
rect 48068 170 48894 272
rect 49008 272 50716 278
rect 49008 264 49822 272
rect 49008 170 49238 264
rect 48068 164 49238 170
rect 47626 148 49238 164
rect 49396 164 49822 264
rect 49936 268 50716 272
rect 49936 164 50336 268
rect 49396 152 50336 164
rect 50494 170 50716 268
rect 50830 170 51494 278
rect 50494 152 51494 170
rect 49396 148 51494 152
rect 46732 142 51494 148
rect 46016 130 51494 142
rect 56544 278 62022 280
rect 56544 272 59422 278
rect 56544 164 56646 272
rect 56760 264 58482 272
rect 56760 258 57996 264
rect 56760 164 57102 258
rect 56544 142 57102 164
rect 57260 256 57996 258
rect 57260 148 57592 256
rect 57706 148 57996 256
rect 58154 164 58482 264
rect 58596 170 59422 272
rect 59536 272 61244 278
rect 59536 264 60350 272
rect 59536 170 59766 264
rect 58596 164 59766 170
rect 58154 148 59766 164
rect 59924 164 60350 264
rect 60464 268 61244 272
rect 60464 164 60864 268
rect 59924 152 60864 164
rect 61022 170 61244 268
rect 61358 170 62022 278
rect 61022 152 62022 170
rect 59924 148 62022 152
rect 57260 142 62022 148
rect 56544 130 62022 142
<< viali >>
rect 10798 7574 10898 7646
rect 11634 7582 11734 7654
rect 12544 7594 12644 7666
rect 13496 7580 13608 7670
rect 14388 7590 14500 7680
rect 15278 7578 15390 7668
rect 16314 7584 16420 7686
rect 17168 7574 17274 7676
rect 18128 7574 18234 7676
rect 18828 7580 18924 7696
rect 19740 7588 19836 7704
rect 20668 7586 20764 7702
rect 21406 7574 21506 7646
rect 22242 7582 22342 7654
rect 23152 7594 23252 7666
rect 24104 7580 24216 7670
rect 24996 7590 25108 7680
rect 25886 7578 25998 7668
rect 26922 7584 27028 7686
rect 27776 7574 27882 7676
rect 28736 7574 28842 7676
rect 29436 7580 29532 7696
rect 30348 7588 30444 7704
rect 31276 7586 31372 7702
rect 31934 7574 32034 7646
rect 32770 7582 32870 7654
rect 33680 7594 33780 7666
rect 34632 7580 34744 7670
rect 35524 7590 35636 7680
rect 36414 7578 36526 7668
rect 37450 7584 37556 7686
rect 38304 7574 38410 7676
rect 39264 7574 39370 7676
rect 39964 7580 40060 7696
rect 40876 7588 40972 7704
rect 41804 7586 41900 7702
rect 42544 7574 42644 7646
rect 43380 7582 43480 7654
rect 44290 7594 44390 7666
rect 45242 7580 45354 7670
rect 46134 7590 46246 7680
rect 47024 7578 47136 7668
rect 48060 7584 48166 7686
rect 48914 7574 49020 7676
rect 49874 7574 49980 7676
rect 50574 7580 50670 7696
rect 51486 7588 51582 7704
rect 52414 7586 52510 7702
rect 53072 7574 53172 7646
rect 53908 7582 54008 7654
rect 54818 7594 54918 7666
rect 55770 7580 55882 7670
rect 56662 7590 56774 7680
rect 57552 7578 57664 7668
rect 58588 7584 58694 7686
rect 59442 7574 59548 7676
rect 60402 7574 60508 7676
rect 61102 7580 61198 7696
rect 62014 7588 62110 7704
rect 62942 7586 63038 7702
rect 10732 7360 10742 7386
rect 10742 7360 10804 7386
rect 14252 7388 14328 7408
rect 10732 7350 10804 7360
rect 10752 7020 10760 7092
rect 10760 7020 10786 7092
rect 11674 7016 11676 7088
rect 11676 7016 11708 7088
rect 11216 6706 11218 6778
rect 11218 6706 11250 6778
rect 12588 7016 12592 7088
rect 12592 7016 12622 7088
rect 12126 6706 12134 6784
rect 12134 6706 12162 6784
rect 10815 5130 10822 5161
rect 10822 5130 11183 5161
rect 11273 5130 11280 5161
rect 11280 5130 11641 5161
rect 11731 5130 11738 5161
rect 11738 5130 12099 5161
rect 12189 5130 12196 5161
rect 12196 5130 12557 5161
rect 10815 5127 11183 5130
rect 11273 5127 11641 5130
rect 11731 5127 12099 5130
rect 12189 5127 12557 5130
rect 14252 7364 14328 7388
rect 19456 7384 19522 7394
rect 16756 7362 16826 7372
rect 13576 7252 13944 7286
rect 14034 7252 14402 7286
rect 14492 7252 14860 7286
rect 14950 7252 15318 7286
rect 13508 7022 13514 7104
rect 13514 7022 13544 7104
rect 14426 7016 14430 7098
rect 14430 7016 14462 7098
rect 13966 6804 13972 6886
rect 13972 6804 14002 6886
rect 15340 7016 15346 7098
rect 15346 7016 15376 7098
rect 14894 6798 14922 6880
rect 14922 6798 14930 6880
rect 16756 7328 16826 7362
rect 16756 7326 16826 7328
rect 16392 7226 16760 7260
rect 16850 7226 17218 7260
rect 17308 7226 17676 7260
rect 17766 7226 18134 7260
rect 16328 7006 16330 7098
rect 16330 7006 16364 7098
rect 16364 7006 16378 7098
rect 17248 7008 17280 7094
rect 17280 7008 17288 7094
rect 16790 6720 16822 6806
rect 16822 6720 16830 6806
rect 18160 7016 18162 7102
rect 18162 7016 18196 7102
rect 18196 7016 18200 7102
rect 17706 6720 17738 6806
rect 17738 6720 17746 6806
rect 19456 7350 19522 7384
rect 18858 7010 18888 7072
rect 18888 7010 18894 7072
rect 19780 7008 19804 7100
rect 19804 7008 19818 7100
rect 19292 6614 19312 6720
rect 19312 6614 19346 6720
rect 19346 6614 19360 6720
rect 20688 7018 20720 7110
rect 20720 7018 20726 7110
rect 20214 6622 20228 6728
rect 20228 6622 20262 6728
rect 20262 6622 20282 6728
rect 18916 5120 19284 5154
rect 19374 5120 19742 5154
rect 19832 5120 20200 5154
rect 20290 5120 20658 5154
rect 21340 7360 21350 7386
rect 21350 7360 21412 7386
rect 24860 7388 24936 7408
rect 21340 7350 21412 7360
rect 21360 7020 21368 7092
rect 21368 7020 21394 7092
rect 22282 7016 22284 7088
rect 22284 7016 22316 7088
rect 21824 6706 21826 6778
rect 21826 6706 21858 6778
rect 23196 7016 23200 7088
rect 23200 7016 23230 7088
rect 22734 6706 22742 6784
rect 22742 6706 22770 6784
rect 21423 5130 21430 5161
rect 21430 5130 21791 5161
rect 21881 5130 21888 5161
rect 21888 5130 22249 5161
rect 22339 5130 22346 5161
rect 22346 5130 22707 5161
rect 22797 5130 22804 5161
rect 22804 5130 23165 5161
rect 21423 5127 21791 5130
rect 21881 5127 22249 5130
rect 22339 5127 22707 5130
rect 22797 5127 23165 5130
rect 24860 7364 24936 7388
rect 30064 7384 30130 7394
rect 27364 7362 27434 7372
rect 24184 7252 24552 7286
rect 24642 7252 25010 7286
rect 25100 7252 25468 7286
rect 25558 7252 25926 7286
rect 24116 7022 24122 7104
rect 24122 7022 24152 7104
rect 25034 7016 25038 7098
rect 25038 7016 25070 7098
rect 24574 6804 24580 6886
rect 24580 6804 24610 6886
rect 25948 7016 25954 7098
rect 25954 7016 25984 7098
rect 25502 6798 25530 6880
rect 25530 6798 25538 6880
rect 27364 7328 27434 7362
rect 27364 7326 27434 7328
rect 27000 7226 27368 7260
rect 27458 7226 27826 7260
rect 27916 7226 28284 7260
rect 28374 7226 28742 7260
rect 26936 7006 26938 7098
rect 26938 7006 26972 7098
rect 26972 7006 26986 7098
rect 27856 7008 27888 7094
rect 27888 7008 27896 7094
rect 27398 6720 27430 6806
rect 27430 6720 27438 6806
rect 28768 7016 28770 7102
rect 28770 7016 28804 7102
rect 28804 7016 28808 7102
rect 28314 6720 28346 6806
rect 28346 6720 28354 6806
rect 30064 7350 30130 7384
rect 29466 7010 29496 7072
rect 29496 7010 29502 7072
rect 30388 7008 30412 7100
rect 30412 7008 30426 7100
rect 29900 6614 29920 6720
rect 29920 6614 29954 6720
rect 29954 6614 29968 6720
rect 31296 7018 31328 7110
rect 31328 7018 31334 7110
rect 30822 6622 30836 6728
rect 30836 6622 30870 6728
rect 30870 6622 30890 6728
rect 29524 5120 29892 5154
rect 29982 5120 30350 5154
rect 30440 5120 30808 5154
rect 30898 5120 31266 5154
rect 31868 7360 31878 7386
rect 31878 7360 31940 7386
rect 35388 7388 35464 7408
rect 31868 7350 31940 7360
rect 31888 7020 31896 7092
rect 31896 7020 31922 7092
rect 32810 7016 32812 7088
rect 32812 7016 32844 7088
rect 32352 6706 32354 6778
rect 32354 6706 32386 6778
rect 33724 7016 33728 7088
rect 33728 7016 33758 7088
rect 33262 6706 33270 6784
rect 33270 6706 33298 6784
rect 31951 5130 31958 5161
rect 31958 5130 32319 5161
rect 32409 5130 32416 5161
rect 32416 5130 32777 5161
rect 32867 5130 32874 5161
rect 32874 5130 33235 5161
rect 33325 5130 33332 5161
rect 33332 5130 33693 5161
rect 31951 5127 32319 5130
rect 32409 5127 32777 5130
rect 32867 5127 33235 5130
rect 33325 5127 33693 5130
rect 35388 7364 35464 7388
rect 40592 7384 40658 7394
rect 37892 7362 37962 7372
rect 34712 7252 35080 7286
rect 35170 7252 35538 7286
rect 35628 7252 35996 7286
rect 36086 7252 36454 7286
rect 34644 7022 34650 7104
rect 34650 7022 34680 7104
rect 35562 7016 35566 7098
rect 35566 7016 35598 7098
rect 35102 6804 35108 6886
rect 35108 6804 35138 6886
rect 36476 7016 36482 7098
rect 36482 7016 36512 7098
rect 36030 6798 36058 6880
rect 36058 6798 36066 6880
rect 37892 7328 37962 7362
rect 37892 7326 37962 7328
rect 37528 7226 37896 7260
rect 37986 7226 38354 7260
rect 38444 7226 38812 7260
rect 38902 7226 39270 7260
rect 37464 7006 37466 7098
rect 37466 7006 37500 7098
rect 37500 7006 37514 7098
rect 38384 7008 38416 7094
rect 38416 7008 38424 7094
rect 37926 6720 37958 6806
rect 37958 6720 37966 6806
rect 39296 7016 39298 7102
rect 39298 7016 39332 7102
rect 39332 7016 39336 7102
rect 38842 6720 38874 6806
rect 38874 6720 38882 6806
rect 40592 7350 40658 7384
rect 39994 7010 40024 7072
rect 40024 7010 40030 7072
rect 40916 7008 40940 7100
rect 40940 7008 40954 7100
rect 40428 6614 40448 6720
rect 40448 6614 40482 6720
rect 40482 6614 40496 6720
rect 41824 7018 41856 7110
rect 41856 7018 41862 7110
rect 41350 6622 41364 6728
rect 41364 6622 41398 6728
rect 41398 6622 41418 6728
rect 40052 5120 40420 5154
rect 40510 5120 40878 5154
rect 40968 5120 41336 5154
rect 41426 5120 41794 5154
rect 42478 7360 42488 7386
rect 42488 7360 42550 7386
rect 45998 7388 46074 7408
rect 42478 7350 42550 7360
rect 42498 7020 42506 7092
rect 42506 7020 42532 7092
rect 43420 7016 43422 7088
rect 43422 7016 43454 7088
rect 42962 6706 42964 6778
rect 42964 6706 42996 6778
rect 44334 7016 44338 7088
rect 44338 7016 44368 7088
rect 43872 6706 43880 6784
rect 43880 6706 43908 6784
rect 42561 5130 42568 5161
rect 42568 5130 42929 5161
rect 43019 5130 43026 5161
rect 43026 5130 43387 5161
rect 43477 5130 43484 5161
rect 43484 5130 43845 5161
rect 43935 5130 43942 5161
rect 43942 5130 44303 5161
rect 42561 5127 42929 5130
rect 43019 5127 43387 5130
rect 43477 5127 43845 5130
rect 43935 5127 44303 5130
rect 45998 7364 46074 7388
rect 51202 7384 51268 7394
rect 48502 7362 48572 7372
rect 45322 7252 45690 7286
rect 45780 7252 46148 7286
rect 46238 7252 46606 7286
rect 46696 7252 47064 7286
rect 45254 7022 45260 7104
rect 45260 7022 45290 7104
rect 46172 7016 46176 7098
rect 46176 7016 46208 7098
rect 45712 6804 45718 6886
rect 45718 6804 45748 6886
rect 47086 7016 47092 7098
rect 47092 7016 47122 7098
rect 46640 6798 46668 6880
rect 46668 6798 46676 6880
rect 48502 7328 48572 7362
rect 48502 7326 48572 7328
rect 48138 7226 48506 7260
rect 48596 7226 48964 7260
rect 49054 7226 49422 7260
rect 49512 7226 49880 7260
rect 48074 7006 48076 7098
rect 48076 7006 48110 7098
rect 48110 7006 48124 7098
rect 48994 7008 49026 7094
rect 49026 7008 49034 7094
rect 48536 6720 48568 6806
rect 48568 6720 48576 6806
rect 49906 7016 49908 7102
rect 49908 7016 49942 7102
rect 49942 7016 49946 7102
rect 49452 6720 49484 6806
rect 49484 6720 49492 6806
rect 51202 7350 51268 7384
rect 50604 7010 50634 7072
rect 50634 7010 50640 7072
rect 51526 7008 51550 7100
rect 51550 7008 51564 7100
rect 51038 6614 51058 6720
rect 51058 6614 51092 6720
rect 51092 6614 51106 6720
rect 52434 7018 52466 7110
rect 52466 7018 52472 7110
rect 51960 6622 51974 6728
rect 51974 6622 52008 6728
rect 52008 6622 52028 6728
rect 50662 5120 51030 5154
rect 51120 5120 51488 5154
rect 51578 5120 51946 5154
rect 52036 5120 52404 5154
rect 53006 7360 53016 7386
rect 53016 7360 53078 7386
rect 56526 7388 56602 7408
rect 53006 7350 53078 7360
rect 53026 7020 53034 7092
rect 53034 7020 53060 7092
rect 53948 7016 53950 7088
rect 53950 7016 53982 7088
rect 53490 6706 53492 6778
rect 53492 6706 53524 6778
rect 54862 7016 54866 7088
rect 54866 7016 54896 7088
rect 54400 6706 54408 6784
rect 54408 6706 54436 6784
rect 53089 5130 53096 5161
rect 53096 5130 53457 5161
rect 53547 5130 53554 5161
rect 53554 5130 53915 5161
rect 54005 5130 54012 5161
rect 54012 5130 54373 5161
rect 54463 5130 54470 5161
rect 54470 5130 54831 5161
rect 53089 5127 53457 5130
rect 53547 5127 53915 5130
rect 54005 5127 54373 5130
rect 54463 5127 54831 5130
rect 56526 7364 56602 7388
rect 61730 7384 61796 7394
rect 59030 7362 59100 7372
rect 55850 7252 56218 7286
rect 56308 7252 56676 7286
rect 56766 7252 57134 7286
rect 57224 7252 57592 7286
rect 55782 7022 55788 7104
rect 55788 7022 55818 7104
rect 56700 7016 56704 7098
rect 56704 7016 56736 7098
rect 56240 6804 56246 6886
rect 56246 6804 56276 6886
rect 57614 7016 57620 7098
rect 57620 7016 57650 7098
rect 57168 6798 57196 6880
rect 57196 6798 57204 6880
rect 59030 7328 59100 7362
rect 59030 7326 59100 7328
rect 58666 7226 59034 7260
rect 59124 7226 59492 7260
rect 59582 7226 59950 7260
rect 60040 7226 60408 7260
rect 58602 7006 58604 7098
rect 58604 7006 58638 7098
rect 58638 7006 58652 7098
rect 59522 7008 59554 7094
rect 59554 7008 59562 7094
rect 59064 6720 59096 6806
rect 59096 6720 59104 6806
rect 60434 7016 60436 7102
rect 60436 7016 60470 7102
rect 60470 7016 60474 7102
rect 59980 6720 60012 6806
rect 60012 6720 60020 6806
rect 61730 7350 61796 7384
rect 61132 7010 61162 7072
rect 61162 7010 61168 7072
rect 62054 7008 62078 7100
rect 62078 7008 62092 7100
rect 61566 6614 61586 6720
rect 61586 6614 61620 6720
rect 61620 6614 61634 6720
rect 62962 7018 62994 7110
rect 62994 7018 63000 7110
rect 62488 6622 62502 6728
rect 62502 6622 62536 6728
rect 62536 6622 62556 6728
rect 61190 5120 61558 5154
rect 61648 5120 62016 5154
rect 62106 5120 62474 5154
rect 62564 5120 62932 5154
rect 12984 4122 13124 4130
rect 12984 4094 13124 4122
rect 12008 4044 12042 4078
rect 13018 4000 13124 4034
rect 13018 3988 13124 4000
rect 13010 3920 13116 3926
rect 13010 3886 13116 3920
rect 18472 4132 18556 4142
rect 18472 4102 18556 4132
rect 19568 4054 19602 4088
rect 18472 4044 18552 4046
rect 18472 4010 18552 4044
rect 18472 4006 18552 4010
rect 18474 3930 18554 3940
rect 18474 3900 18554 3930
rect 23592 4122 23732 4130
rect 23592 4094 23732 4122
rect 22616 4044 22650 4078
rect 23626 4000 23732 4034
rect 23626 3988 23732 4000
rect 23618 3920 23724 3926
rect 23618 3886 23724 3920
rect 29080 4132 29164 4142
rect 29080 4102 29164 4132
rect 30176 4054 30210 4088
rect 29080 4044 29160 4046
rect 29080 4010 29160 4044
rect 29080 4006 29160 4010
rect 29082 3930 29162 3940
rect 29082 3900 29162 3930
rect 34120 4122 34260 4130
rect 34120 4094 34260 4122
rect 33144 4044 33178 4078
rect 34154 4000 34260 4034
rect 34154 3988 34260 4000
rect 34146 3920 34252 3926
rect 34146 3886 34252 3920
rect 39608 4132 39692 4142
rect 39608 4102 39692 4132
rect 40704 4054 40738 4088
rect 39608 4044 39688 4046
rect 39608 4010 39688 4044
rect 39608 4006 39688 4010
rect 39610 3930 39690 3940
rect 39610 3900 39690 3930
rect 44730 4122 44870 4130
rect 44730 4094 44870 4122
rect 43754 4044 43788 4078
rect 44764 4000 44870 4034
rect 44764 3988 44870 4000
rect 44756 3920 44862 3926
rect 44756 3886 44862 3920
rect 50218 4132 50302 4142
rect 50218 4102 50302 4132
rect 51314 4054 51348 4088
rect 50218 4044 50298 4046
rect 50218 4010 50298 4044
rect 50218 4006 50298 4010
rect 50220 3930 50300 3940
rect 50220 3900 50300 3930
rect 55258 4122 55398 4130
rect 55258 4094 55398 4122
rect 54282 4044 54316 4078
rect 55292 4000 55398 4034
rect 55292 3988 55398 4000
rect 55284 3920 55390 3926
rect 55284 3886 55390 3920
rect 60746 4132 60830 4142
rect 60746 4102 60830 4132
rect 61842 4054 61876 4088
rect 60746 4044 60826 4046
rect 60746 4010 60826 4044
rect 60746 4006 60826 4010
rect 60748 3930 60828 3940
rect 60748 3900 60828 3930
rect 13010 3880 13116 3886
rect 23618 3880 23724 3886
rect 34146 3880 34252 3886
rect 44756 3880 44862 3886
rect 55284 3880 55390 3886
rect 14422 2862 14429 2958
rect 14429 2862 14463 2958
rect 14463 2862 14470 2958
rect 15338 2854 15345 2950
rect 15345 2854 15379 2950
rect 15379 2854 15386 2950
rect 14854 2646 14887 2756
rect 14887 2646 14921 2756
rect 14921 2646 14924 2756
rect 16256 2866 16261 2962
rect 16261 2866 16295 2962
rect 16295 2866 16304 2962
rect 15778 2658 15803 2768
rect 15803 2658 15837 2768
rect 15837 2658 15848 2768
rect 17164 2874 17177 2970
rect 17177 2874 17211 2970
rect 17211 2874 17212 2970
rect 16696 2670 16719 2780
rect 16719 2670 16753 2780
rect 16753 2670 16766 2780
rect 18070 2868 18093 2964
rect 18093 2868 18118 2964
rect 17620 2670 17635 2780
rect 17635 2670 17669 2780
rect 17669 2670 17690 2780
rect 19002 2868 19009 2964
rect 19009 2868 19043 2964
rect 19043 2868 19050 2964
rect 18544 2658 18551 2768
rect 18551 2658 18585 2768
rect 18585 2658 18614 2768
rect 19440 2676 19467 2786
rect 19467 2676 19501 2786
rect 19501 2676 19510 2786
rect 14491 581 14859 615
rect 14949 581 15317 615
rect 15407 581 15775 615
rect 15865 581 16233 615
rect 16323 581 16691 615
rect 16781 581 17149 615
rect 17239 581 17607 615
rect 17697 581 18065 615
rect 18155 581 18523 615
rect 18613 581 18981 615
rect 19071 581 19439 615
rect 18344 479 18446 504
rect 25030 2862 25037 2958
rect 25037 2862 25071 2958
rect 25071 2862 25078 2958
rect 25946 2854 25953 2950
rect 25953 2854 25987 2950
rect 25987 2854 25994 2950
rect 25462 2646 25495 2756
rect 25495 2646 25529 2756
rect 25529 2646 25532 2756
rect 26864 2866 26869 2962
rect 26869 2866 26903 2962
rect 26903 2866 26912 2962
rect 26386 2658 26411 2768
rect 26411 2658 26445 2768
rect 26445 2658 26456 2768
rect 27772 2874 27785 2970
rect 27785 2874 27819 2970
rect 27819 2874 27820 2970
rect 27304 2670 27327 2780
rect 27327 2670 27361 2780
rect 27361 2670 27374 2780
rect 28678 2868 28701 2964
rect 28701 2868 28726 2964
rect 28228 2670 28243 2780
rect 28243 2670 28277 2780
rect 28277 2670 28298 2780
rect 29610 2868 29617 2964
rect 29617 2868 29651 2964
rect 29651 2868 29658 2964
rect 29152 2658 29159 2768
rect 29159 2658 29193 2768
rect 29193 2658 29222 2768
rect 30048 2676 30075 2786
rect 30075 2676 30109 2786
rect 30109 2676 30118 2786
rect 25099 581 25467 615
rect 25557 581 25925 615
rect 26015 581 26383 615
rect 26473 581 26841 615
rect 26931 581 27299 615
rect 27389 581 27757 615
rect 27847 581 28215 615
rect 28305 581 28673 615
rect 28763 581 29131 615
rect 29221 581 29589 615
rect 29679 581 30047 615
rect 28952 479 29054 504
rect 35558 2862 35565 2958
rect 35565 2862 35599 2958
rect 35599 2862 35606 2958
rect 36474 2854 36481 2950
rect 36481 2854 36515 2950
rect 36515 2854 36522 2950
rect 35990 2646 36023 2756
rect 36023 2646 36057 2756
rect 36057 2646 36060 2756
rect 37392 2866 37397 2962
rect 37397 2866 37431 2962
rect 37431 2866 37440 2962
rect 36914 2658 36939 2768
rect 36939 2658 36973 2768
rect 36973 2658 36984 2768
rect 38300 2874 38313 2970
rect 38313 2874 38347 2970
rect 38347 2874 38348 2970
rect 37832 2670 37855 2780
rect 37855 2670 37889 2780
rect 37889 2670 37902 2780
rect 39206 2868 39229 2964
rect 39229 2868 39254 2964
rect 38756 2670 38771 2780
rect 38771 2670 38805 2780
rect 38805 2670 38826 2780
rect 40138 2868 40145 2964
rect 40145 2868 40179 2964
rect 40179 2868 40186 2964
rect 39680 2658 39687 2768
rect 39687 2658 39721 2768
rect 39721 2658 39750 2768
rect 40576 2676 40603 2786
rect 40603 2676 40637 2786
rect 40637 2676 40646 2786
rect 35627 581 35995 615
rect 36085 581 36453 615
rect 36543 581 36911 615
rect 37001 581 37369 615
rect 37459 581 37827 615
rect 37917 581 38285 615
rect 38375 581 38743 615
rect 38833 581 39201 615
rect 39291 581 39659 615
rect 39749 581 40117 615
rect 40207 581 40575 615
rect 39480 479 39582 504
rect 46168 2862 46175 2958
rect 46175 2862 46209 2958
rect 46209 2862 46216 2958
rect 47084 2854 47091 2950
rect 47091 2854 47125 2950
rect 47125 2854 47132 2950
rect 46600 2646 46633 2756
rect 46633 2646 46667 2756
rect 46667 2646 46670 2756
rect 48002 2866 48007 2962
rect 48007 2866 48041 2962
rect 48041 2866 48050 2962
rect 47524 2658 47549 2768
rect 47549 2658 47583 2768
rect 47583 2658 47594 2768
rect 48910 2874 48923 2970
rect 48923 2874 48957 2970
rect 48957 2874 48958 2970
rect 48442 2670 48465 2780
rect 48465 2670 48499 2780
rect 48499 2670 48512 2780
rect 49816 2868 49839 2964
rect 49839 2868 49864 2964
rect 49366 2670 49381 2780
rect 49381 2670 49415 2780
rect 49415 2670 49436 2780
rect 50748 2868 50755 2964
rect 50755 2868 50789 2964
rect 50789 2868 50796 2964
rect 50290 2658 50297 2768
rect 50297 2658 50331 2768
rect 50331 2658 50360 2768
rect 51186 2676 51213 2786
rect 51213 2676 51247 2786
rect 51247 2676 51256 2786
rect 46237 581 46605 615
rect 46695 581 47063 615
rect 47153 581 47521 615
rect 47611 581 47979 615
rect 48069 581 48437 615
rect 48527 581 48895 615
rect 48985 581 49353 615
rect 49443 581 49811 615
rect 49901 581 50269 615
rect 50359 581 50727 615
rect 50817 581 51185 615
rect 50090 479 50192 504
rect 56696 2862 56703 2958
rect 56703 2862 56737 2958
rect 56737 2862 56744 2958
rect 57612 2854 57619 2950
rect 57619 2854 57653 2950
rect 57653 2854 57660 2950
rect 57128 2646 57161 2756
rect 57161 2646 57195 2756
rect 57195 2646 57198 2756
rect 58530 2866 58535 2962
rect 58535 2866 58569 2962
rect 58569 2866 58578 2962
rect 58052 2658 58077 2768
rect 58077 2658 58111 2768
rect 58111 2658 58122 2768
rect 59438 2874 59451 2970
rect 59451 2874 59485 2970
rect 59485 2874 59486 2970
rect 58970 2670 58993 2780
rect 58993 2670 59027 2780
rect 59027 2670 59040 2780
rect 60344 2868 60367 2964
rect 60367 2868 60392 2964
rect 59894 2670 59909 2780
rect 59909 2670 59943 2780
rect 59943 2670 59964 2780
rect 61276 2868 61283 2964
rect 61283 2868 61317 2964
rect 61317 2868 61324 2964
rect 60818 2658 60825 2768
rect 60825 2658 60859 2768
rect 60859 2658 60888 2768
rect 61714 2676 61741 2786
rect 61741 2676 61775 2786
rect 61775 2676 61784 2786
rect 56765 581 57133 615
rect 57223 581 57591 615
rect 57681 581 58049 615
rect 58139 581 58507 615
rect 58597 581 58965 615
rect 59055 581 59423 615
rect 59513 581 59881 615
rect 59971 581 60339 615
rect 60429 581 60797 615
rect 60887 581 61255 615
rect 61345 581 61713 615
rect 60618 479 60720 504
rect 18344 470 18446 479
rect 28952 470 29054 479
rect 39480 470 39582 479
rect 50090 470 50192 479
rect 60618 470 60720 479
rect 14372 164 14486 272
rect 15318 148 15432 256
rect 16208 164 16322 272
rect 17148 170 17262 278
rect 18076 164 18190 272
rect 18970 170 19084 278
rect 24980 164 25094 272
rect 25926 148 26040 256
rect 26816 164 26930 272
rect 27756 170 27870 278
rect 28684 164 28798 272
rect 29578 170 29692 278
rect 35508 164 35622 272
rect 36454 148 36568 256
rect 37344 164 37458 272
rect 38284 170 38398 278
rect 39212 164 39326 272
rect 40106 170 40220 278
rect 46118 164 46232 272
rect 47064 148 47178 256
rect 47954 164 48068 272
rect 48894 170 49008 278
rect 49822 164 49936 272
rect 50716 170 50830 278
rect 56646 164 56760 272
rect 57592 148 57706 256
rect 58482 164 58596 272
rect 59422 170 59536 278
rect 60350 164 60464 272
rect 61244 170 61358 278
<< metal1 >>
rect 3057 8000 11488 8470
rect 3057 7704 63264 8000
rect 3057 7696 19740 7704
rect 3057 7686 16320 7696
rect 16374 7686 18828 7696
rect 3057 7680 16314 7686
rect 3057 7670 14388 7680
rect 3057 7666 13496 7670
rect 3057 7654 12544 7666
rect 3057 7646 11634 7654
rect 3057 7574 10798 7646
rect 10898 7582 11634 7646
rect 11734 7594 12544 7654
rect 12644 7594 13496 7666
rect 11734 7582 13496 7594
rect 10898 7580 13496 7582
rect 13608 7590 14388 7670
rect 14500 7668 16314 7680
rect 14500 7590 15278 7668
rect 13608 7580 15278 7590
rect 10898 7578 15278 7580
rect 15390 7584 16314 7668
rect 16420 7676 18828 7686
rect 16420 7584 17168 7676
rect 15390 7578 17168 7584
rect 10898 7574 17168 7578
rect 17274 7574 18128 7676
rect 18234 7580 18828 7676
rect 18924 7588 19740 7696
rect 19836 7702 30348 7704
rect 19836 7588 20668 7702
rect 18924 7586 20668 7588
rect 20764 7696 30348 7702
rect 20764 7686 26928 7696
rect 26982 7686 29436 7696
rect 20764 7680 26922 7686
rect 20764 7670 24996 7680
rect 20764 7666 24104 7670
rect 20764 7654 23152 7666
rect 20764 7646 22242 7654
rect 20764 7586 21406 7646
rect 18924 7580 21406 7586
rect 18234 7574 21406 7580
rect 21506 7582 22242 7646
rect 22342 7594 23152 7654
rect 23252 7594 24104 7666
rect 22342 7582 24104 7594
rect 21506 7580 24104 7582
rect 24216 7590 24996 7670
rect 25108 7668 26922 7680
rect 25108 7590 25886 7668
rect 24216 7580 25886 7590
rect 21506 7578 25886 7580
rect 25998 7584 26922 7668
rect 27028 7676 29436 7686
rect 27028 7584 27776 7676
rect 25998 7578 27776 7584
rect 21506 7574 27776 7578
rect 27882 7574 28736 7676
rect 28842 7580 29436 7676
rect 29532 7588 30348 7696
rect 30444 7702 40876 7704
rect 30444 7588 31276 7702
rect 29532 7586 31276 7588
rect 31372 7696 40876 7702
rect 31372 7686 37456 7696
rect 37510 7686 39964 7696
rect 31372 7680 37450 7686
rect 31372 7670 35524 7680
rect 31372 7666 34632 7670
rect 31372 7654 33680 7666
rect 31372 7646 32770 7654
rect 31372 7586 31934 7646
rect 29532 7580 31934 7586
rect 28842 7574 31934 7580
rect 32034 7582 32770 7646
rect 32870 7594 33680 7654
rect 33780 7594 34632 7666
rect 32870 7582 34632 7594
rect 32034 7580 34632 7582
rect 34744 7590 35524 7670
rect 35636 7668 37450 7680
rect 35636 7590 36414 7668
rect 34744 7580 36414 7590
rect 32034 7578 36414 7580
rect 36526 7584 37450 7668
rect 37556 7676 39964 7686
rect 37556 7584 38304 7676
rect 36526 7578 38304 7584
rect 32034 7574 38304 7578
rect 38410 7574 39264 7676
rect 39370 7580 39964 7676
rect 40060 7588 40876 7696
rect 40972 7702 51486 7704
rect 40972 7588 41804 7702
rect 40060 7586 41804 7588
rect 41900 7696 51486 7702
rect 41900 7686 48066 7696
rect 48120 7686 50574 7696
rect 41900 7680 48060 7686
rect 41900 7670 46134 7680
rect 41900 7666 45242 7670
rect 41900 7654 44290 7666
rect 41900 7646 43380 7654
rect 41900 7586 42544 7646
rect 40060 7580 42544 7586
rect 39370 7574 42544 7580
rect 42644 7582 43380 7646
rect 43480 7594 44290 7654
rect 44390 7594 45242 7666
rect 43480 7582 45242 7594
rect 42644 7580 45242 7582
rect 45354 7590 46134 7670
rect 46246 7668 48060 7680
rect 46246 7590 47024 7668
rect 45354 7580 47024 7590
rect 42644 7578 47024 7580
rect 47136 7584 48060 7668
rect 48166 7676 50574 7686
rect 48166 7584 48914 7676
rect 47136 7578 48914 7584
rect 42644 7574 48914 7578
rect 49020 7574 49874 7676
rect 49980 7580 50574 7676
rect 50670 7588 51486 7696
rect 51582 7702 62014 7704
rect 51582 7588 52414 7702
rect 50670 7586 52414 7588
rect 52510 7696 62014 7702
rect 52510 7686 58594 7696
rect 58648 7686 61102 7696
rect 52510 7680 58588 7686
rect 52510 7670 56662 7680
rect 52510 7666 55770 7670
rect 52510 7654 54818 7666
rect 52510 7646 53908 7654
rect 52510 7586 53072 7646
rect 50670 7580 53072 7586
rect 49980 7574 53072 7580
rect 53172 7582 53908 7646
rect 54008 7594 54818 7654
rect 54918 7594 55770 7666
rect 54008 7582 55770 7594
rect 53172 7580 55770 7582
rect 55882 7590 56662 7670
rect 56774 7668 58588 7680
rect 56774 7590 57552 7668
rect 55882 7580 57552 7590
rect 53172 7578 57552 7580
rect 57664 7584 58588 7668
rect 58694 7676 61102 7686
rect 58694 7584 59442 7676
rect 57664 7578 59442 7584
rect 53172 7574 59442 7578
rect 59548 7574 60402 7676
rect 60508 7580 61102 7676
rect 61198 7588 62014 7696
rect 62110 7702 63264 7704
rect 62110 7588 62942 7702
rect 61198 7586 62942 7588
rect 63038 7586 63264 7702
rect 61198 7580 63264 7586
rect 60508 7574 63264 7580
rect 3057 7523 63264 7574
rect 10548 7510 63264 7523
rect 10704 7386 10822 7510
rect 10704 7350 10732 7386
rect 10804 7350 10822 7386
rect 10704 7102 10822 7350
rect 14238 7408 14344 7510
rect 14238 7364 14252 7408
rect 14328 7364 14344 7408
rect 14238 7346 14344 7364
rect 16736 7372 16862 7510
rect 15722 7314 16011 7351
rect 16736 7326 16756 7372
rect 16826 7326 16862 7372
rect 16736 7318 16862 7326
rect 13536 7304 16344 7314
rect 13536 7286 15765 7304
rect 13536 7252 13576 7286
rect 13944 7252 14034 7286
rect 14402 7252 14492 7286
rect 14860 7252 14950 7286
rect 15318 7252 15765 7286
rect 13536 7220 15765 7252
rect 15514 7194 15765 7220
rect 15722 7185 15765 7194
rect 15972 7278 16344 7304
rect 15972 7260 18196 7278
rect 15972 7226 16392 7260
rect 16760 7226 16850 7260
rect 17218 7226 17308 7260
rect 17676 7226 17766 7260
rect 18134 7226 18196 7260
rect 15972 7194 18196 7226
rect 15972 7185 16011 7194
rect 15722 7142 16011 7185
rect 18836 7122 18918 7510
rect 19442 7500 20990 7510
rect 19442 7394 19540 7500
rect 19442 7350 19456 7394
rect 19522 7350 19540 7394
rect 19442 7336 19540 7350
rect 21312 7386 21430 7510
rect 21312 7350 21340 7386
rect 21412 7350 21430 7386
rect 13470 7104 15422 7118
rect 12094 7102 12384 7104
rect 10704 7092 12658 7102
rect 10704 7020 10752 7092
rect 10786 7088 12658 7092
rect 10786 7020 11674 7088
rect 10704 7016 11674 7020
rect 11708 7016 12588 7088
rect 12622 7016 12658 7088
rect 10704 7014 12658 7016
rect 10704 7006 12196 7014
rect 12280 7006 12658 7014
rect 13470 7094 13508 7104
rect 13544 7098 15422 7104
rect 13544 7094 14426 7098
rect 13470 7002 13500 7094
rect 13606 7016 14426 7094
rect 14462 7016 15340 7098
rect 15376 7016 15422 7098
rect 13606 7002 15422 7016
rect 13470 6988 15422 7002
rect 16290 7102 18252 7118
rect 16290 7098 18160 7102
rect 16290 7088 16328 7098
rect 16378 7094 18160 7098
rect 16290 6998 16318 7088
rect 16378 7008 17248 7094
rect 17288 7016 18160 7094
rect 18200 7016 18252 7102
rect 17288 7008 18252 7016
rect 16378 7006 18252 7008
rect 16372 6998 18252 7006
rect 16290 6986 18252 6998
rect 18832 7110 20744 7122
rect 18832 7100 20688 7110
rect 18832 7072 19780 7100
rect 18832 7010 18858 7072
rect 18894 7010 19780 7072
rect 18832 7008 19780 7010
rect 19818 7018 20688 7100
rect 20726 7018 20744 7110
rect 19818 7008 20744 7018
rect 18832 6970 20744 7008
rect 21312 7102 21430 7350
rect 24846 7408 24952 7510
rect 24846 7364 24860 7408
rect 24936 7364 24952 7408
rect 24846 7346 24952 7364
rect 27344 7372 27470 7510
rect 26332 7314 26621 7346
rect 27344 7326 27364 7372
rect 27434 7326 27470 7372
rect 27344 7318 27470 7326
rect 24144 7299 26952 7314
rect 24144 7286 26375 7299
rect 24144 7252 24184 7286
rect 24552 7252 24642 7286
rect 25010 7252 25100 7286
rect 25468 7252 25558 7286
rect 25926 7252 26375 7286
rect 24144 7220 26375 7252
rect 26122 7194 26375 7220
rect 26332 7180 26375 7194
rect 26582 7278 26952 7299
rect 26582 7260 28804 7278
rect 26582 7226 27000 7260
rect 27368 7226 27458 7260
rect 27826 7226 27916 7260
rect 28284 7226 28374 7260
rect 28742 7226 28804 7260
rect 26582 7194 28804 7226
rect 26582 7180 26621 7194
rect 26332 7137 26621 7180
rect 29444 7122 29526 7510
rect 30050 7500 31598 7510
rect 30050 7394 30148 7500
rect 30050 7350 30064 7394
rect 30130 7350 30148 7394
rect 30050 7336 30148 7350
rect 31840 7386 31958 7510
rect 31840 7350 31868 7386
rect 31940 7350 31958 7386
rect 24078 7104 26030 7118
rect 22702 7102 22992 7104
rect 21312 7092 23266 7102
rect 21312 7020 21360 7092
rect 21394 7088 23266 7092
rect 21394 7020 22282 7088
rect 21312 7016 22282 7020
rect 22316 7016 23196 7088
rect 23230 7016 23266 7088
rect 21312 7014 23266 7016
rect 21312 7006 22804 7014
rect 22888 7006 23266 7014
rect 24078 7094 24116 7104
rect 24152 7098 26030 7104
rect 24152 7094 25034 7098
rect 24078 7002 24108 7094
rect 24214 7016 25034 7094
rect 25070 7016 25948 7098
rect 25984 7016 26030 7098
rect 24214 7002 26030 7016
rect 24078 6988 26030 7002
rect 26898 7102 28860 7118
rect 26898 7098 28768 7102
rect 26898 7088 26936 7098
rect 26986 7094 28768 7098
rect 26898 6998 26926 7088
rect 26986 7008 27856 7094
rect 27896 7016 28768 7094
rect 28808 7016 28860 7102
rect 27896 7008 28860 7016
rect 26986 7006 28860 7008
rect 26980 6998 28860 7006
rect 26898 6986 28860 6998
rect 29440 7110 31352 7122
rect 29440 7100 31296 7110
rect 29440 7072 30388 7100
rect 29440 7010 29466 7072
rect 29502 7010 30388 7072
rect 29440 7008 30388 7010
rect 30426 7018 31296 7100
rect 31334 7018 31352 7110
rect 30426 7008 31352 7018
rect 29440 6970 31352 7008
rect 31840 7102 31958 7350
rect 35374 7408 35480 7510
rect 35374 7364 35388 7408
rect 35464 7364 35480 7408
rect 35374 7346 35480 7364
rect 37872 7372 37998 7510
rect 36861 7314 37150 7346
rect 37872 7326 37892 7372
rect 37962 7326 37998 7372
rect 37872 7318 37998 7326
rect 34672 7299 37480 7314
rect 34672 7286 36904 7299
rect 34672 7252 34712 7286
rect 35080 7252 35170 7286
rect 35538 7252 35628 7286
rect 35996 7252 36086 7286
rect 36454 7252 36904 7286
rect 34672 7220 36904 7252
rect 36650 7194 36904 7220
rect 36861 7180 36904 7194
rect 37111 7278 37480 7299
rect 37111 7260 39332 7278
rect 37111 7226 37528 7260
rect 37896 7226 37986 7260
rect 38354 7226 38444 7260
rect 38812 7226 38902 7260
rect 39270 7226 39332 7260
rect 37111 7194 39332 7226
rect 37111 7180 37150 7194
rect 36861 7137 37150 7180
rect 39972 7122 40054 7510
rect 40578 7500 42126 7510
rect 40578 7394 40676 7500
rect 40578 7350 40592 7394
rect 40658 7350 40676 7394
rect 40578 7336 40676 7350
rect 42450 7386 42568 7510
rect 42450 7350 42478 7386
rect 42550 7350 42568 7386
rect 34606 7104 36558 7118
rect 33230 7102 33520 7104
rect 31840 7092 33794 7102
rect 31840 7020 31888 7092
rect 31922 7088 33794 7092
rect 31922 7020 32810 7088
rect 31840 7016 32810 7020
rect 32844 7016 33724 7088
rect 33758 7016 33794 7088
rect 31840 7014 33794 7016
rect 31840 7006 33332 7014
rect 33416 7006 33794 7014
rect 34606 7094 34644 7104
rect 34680 7098 36558 7104
rect 34680 7094 35562 7098
rect 34606 7002 34636 7094
rect 34742 7016 35562 7094
rect 35598 7016 36476 7098
rect 36512 7016 36558 7098
rect 34742 7002 36558 7016
rect 34606 6988 36558 7002
rect 37426 7102 39388 7118
rect 37426 7098 39296 7102
rect 37426 7088 37464 7098
rect 37514 7094 39296 7098
rect 37426 6998 37454 7088
rect 37514 7008 38384 7094
rect 38424 7016 39296 7094
rect 39336 7016 39388 7102
rect 38424 7008 39388 7016
rect 37514 7006 39388 7008
rect 37508 6998 39388 7006
rect 37426 6986 39388 6998
rect 39968 7110 41880 7122
rect 39968 7100 41824 7110
rect 39968 7072 40916 7100
rect 39968 7010 39994 7072
rect 40030 7010 40916 7072
rect 39968 7008 40916 7010
rect 40954 7018 41824 7100
rect 41862 7018 41880 7110
rect 40954 7008 41880 7018
rect 39968 6970 41880 7008
rect 42450 7102 42568 7350
rect 45984 7408 46090 7510
rect 45984 7364 45998 7408
rect 46074 7364 46090 7408
rect 45984 7346 46090 7364
rect 48482 7372 48608 7510
rect 47444 7314 47733 7346
rect 48482 7326 48502 7372
rect 48572 7326 48608 7372
rect 48482 7318 48608 7326
rect 45282 7299 48090 7314
rect 45282 7286 47487 7299
rect 45282 7252 45322 7286
rect 45690 7252 45780 7286
rect 46148 7252 46238 7286
rect 46606 7252 46696 7286
rect 47064 7252 47487 7286
rect 45282 7220 47487 7252
rect 47260 7194 47487 7220
rect 47444 7180 47487 7194
rect 47694 7278 48090 7299
rect 47694 7260 49942 7278
rect 47694 7226 48138 7260
rect 48506 7226 48596 7260
rect 48964 7226 49054 7260
rect 49422 7226 49512 7260
rect 49880 7226 49942 7260
rect 47694 7194 49942 7226
rect 47694 7180 47733 7194
rect 47444 7137 47733 7180
rect 50582 7122 50664 7510
rect 51188 7500 52736 7510
rect 51188 7394 51286 7500
rect 51188 7350 51202 7394
rect 51268 7350 51286 7394
rect 51188 7336 51286 7350
rect 52978 7386 53096 7510
rect 52978 7350 53006 7386
rect 53078 7350 53096 7386
rect 45216 7104 47168 7118
rect 43840 7102 44130 7104
rect 42450 7092 44404 7102
rect 42450 7020 42498 7092
rect 42532 7088 44404 7092
rect 42532 7020 43420 7088
rect 42450 7016 43420 7020
rect 43454 7016 44334 7088
rect 44368 7016 44404 7088
rect 42450 7014 44404 7016
rect 42450 7006 43942 7014
rect 44026 7006 44404 7014
rect 45216 7094 45254 7104
rect 45290 7098 47168 7104
rect 45290 7094 46172 7098
rect 45216 7002 45246 7094
rect 45352 7016 46172 7094
rect 46208 7016 47086 7098
rect 47122 7016 47168 7098
rect 45352 7002 47168 7016
rect 45216 6988 47168 7002
rect 48036 7102 49998 7118
rect 48036 7098 49906 7102
rect 48036 7088 48074 7098
rect 48124 7094 49906 7098
rect 48036 6998 48064 7088
rect 48124 7008 48994 7094
rect 49034 7016 49906 7094
rect 49946 7016 49998 7102
rect 49034 7008 49998 7016
rect 48124 7006 49998 7008
rect 48118 6998 49998 7006
rect 48036 6986 49998 6998
rect 50578 7110 52490 7122
rect 50578 7100 52434 7110
rect 50578 7072 51526 7100
rect 50578 7010 50604 7072
rect 50640 7010 51526 7072
rect 50578 7008 51526 7010
rect 51564 7018 52434 7100
rect 52472 7018 52490 7110
rect 51564 7008 52490 7018
rect 50578 6970 52490 7008
rect 52978 7102 53096 7350
rect 56512 7408 56618 7510
rect 56512 7364 56526 7408
rect 56602 7364 56618 7408
rect 56512 7346 56618 7364
rect 59010 7372 59136 7510
rect 58014 7328 58303 7360
rect 58002 7314 58317 7328
rect 59010 7326 59030 7372
rect 59100 7326 59136 7372
rect 59010 7318 59136 7326
rect 55810 7313 58618 7314
rect 55810 7286 58057 7313
rect 55810 7252 55850 7286
rect 56218 7252 56308 7286
rect 56676 7252 56766 7286
rect 57134 7252 57224 7286
rect 57592 7252 58057 7286
rect 55810 7220 58057 7252
rect 57788 7194 58057 7220
rect 58264 7278 58618 7313
rect 58264 7260 60470 7278
rect 58264 7226 58666 7260
rect 59034 7226 59124 7260
rect 59492 7226 59582 7260
rect 59950 7226 60040 7260
rect 60408 7226 60470 7260
rect 58264 7194 60470 7226
rect 58014 7151 58303 7194
rect 61110 7122 61192 7510
rect 61716 7500 63264 7510
rect 61716 7394 61814 7500
rect 61716 7350 61730 7394
rect 61796 7350 61814 7394
rect 61716 7336 61814 7350
rect 55744 7104 57696 7118
rect 54368 7102 54658 7104
rect 52978 7092 54932 7102
rect 52978 7020 53026 7092
rect 53060 7088 54932 7092
rect 53060 7020 53948 7088
rect 52978 7016 53948 7020
rect 53982 7016 54862 7088
rect 54896 7016 54932 7088
rect 52978 7014 54932 7016
rect 52978 7006 54470 7014
rect 54554 7006 54932 7014
rect 55744 7094 55782 7104
rect 55818 7098 57696 7104
rect 55818 7094 56700 7098
rect 55744 7002 55774 7094
rect 55880 7016 56700 7094
rect 56736 7016 57614 7098
rect 57650 7016 57696 7098
rect 55880 7002 57696 7016
rect 55744 6988 57696 7002
rect 58564 7102 60526 7118
rect 58564 7098 60434 7102
rect 58564 7088 58602 7098
rect 58652 7094 60434 7098
rect 58564 6998 58592 7088
rect 58652 7008 59522 7094
rect 59562 7016 60434 7094
rect 60474 7016 60526 7102
rect 59562 7008 60526 7016
rect 58652 7006 60526 7008
rect 58646 6998 60526 7006
rect 58564 6986 60526 6998
rect 61106 7110 63018 7122
rect 61106 7100 62962 7110
rect 61106 7072 62054 7100
rect 61106 7010 61132 7072
rect 61168 7010 62054 7072
rect 61106 7008 62054 7010
rect 62092 7018 62962 7100
rect 63000 7018 63018 7110
rect 62092 7008 63018 7018
rect 61106 6970 63018 7008
rect 13952 6894 14944 6900
rect 24560 6894 25552 6900
rect 35088 6894 36080 6900
rect 45698 6894 46690 6900
rect 56226 6894 57218 6900
rect 13926 6886 14944 6894
rect 11160 6784 12196 6806
rect 11160 6778 12126 6784
rect 11160 6706 11216 6778
rect 11250 6706 12126 6778
rect 12162 6706 12196 6784
rect 11160 6684 12196 6706
rect 13926 6804 13966 6886
rect 14002 6880 14944 6886
rect 14002 6804 14894 6880
rect 13926 6798 14894 6804
rect 14930 6798 14944 6880
rect 24534 6886 25552 6894
rect 13926 6766 14944 6798
rect 16758 6806 17784 6834
rect 12058 5178 12190 6684
rect 10754 5161 12608 5178
rect 10754 5127 10815 5161
rect 11183 5127 11273 5161
rect 11641 5127 11731 5161
rect 12099 5127 12189 5161
rect 12557 5127 12608 5161
rect 10754 5090 12608 5127
rect 12058 4910 12190 5090
rect 13926 4910 14056 6766
rect 16758 6720 16790 6806
rect 16830 6720 17706 6806
rect 17746 6720 17784 6806
rect 21768 6784 22804 6806
rect 21768 6778 22734 6784
rect 19272 6760 20302 6764
rect 16758 6702 17784 6720
rect 19262 6728 20302 6760
rect 19262 6720 20214 6728
rect 17648 4914 17780 6702
rect 19262 6614 19292 6720
rect 19360 6622 20214 6720
rect 20282 6622 20302 6728
rect 21768 6706 21824 6778
rect 21858 6706 22734 6778
rect 22770 6706 22804 6784
rect 21768 6684 22804 6706
rect 24534 6804 24574 6886
rect 24610 6880 25552 6886
rect 24610 6804 25502 6880
rect 24534 6798 25502 6804
rect 25538 6798 25552 6880
rect 35062 6886 36080 6894
rect 24534 6766 25552 6798
rect 27366 6806 28392 6834
rect 19360 6614 20302 6622
rect 19262 6584 20302 6614
rect 19262 5178 19384 6584
rect 22666 5178 22798 6684
rect 18868 5154 20704 5178
rect 18868 5120 18916 5154
rect 19284 5120 19374 5154
rect 19742 5120 19832 5154
rect 20200 5120 20290 5154
rect 20658 5120 20704 5154
rect 18868 5102 20704 5120
rect 21362 5161 23216 5178
rect 21362 5127 21423 5161
rect 21791 5127 21881 5161
rect 22249 5127 22339 5161
rect 22707 5127 22797 5161
rect 23165 5127 23216 5161
rect 19262 4970 19384 5102
rect 21362 5090 23216 5127
rect 19262 4914 19382 4970
rect 12058 4878 14056 4910
rect 12058 4780 14062 4878
rect 17644 4869 19382 4914
rect 17644 4830 18476 4869
rect 12958 4636 13176 4780
rect 12958 4499 12996 4636
rect 13134 4499 13176 4636
rect 12958 4130 13176 4499
rect 10854 4090 12060 4096
rect 10854 4033 10871 4090
rect 11557 4078 12060 4090
rect 12958 4094 12984 4130
rect 13124 4094 13176 4130
rect 12958 4080 13176 4094
rect 18454 4772 18476 4830
rect 18551 4830 19382 4869
rect 22666 4910 22798 5090
rect 24534 4910 24664 6766
rect 27366 6720 27398 6806
rect 27438 6720 28314 6806
rect 28354 6720 28392 6806
rect 32296 6784 33332 6806
rect 32296 6778 33262 6784
rect 29880 6760 30910 6764
rect 27366 6702 28392 6720
rect 29870 6728 30910 6760
rect 29870 6720 30822 6728
rect 28256 4914 28388 6702
rect 29870 6614 29900 6720
rect 29968 6622 30822 6720
rect 30890 6622 30910 6728
rect 32296 6706 32352 6778
rect 32386 6706 33262 6778
rect 33298 6706 33332 6784
rect 32296 6684 33332 6706
rect 35062 6804 35102 6886
rect 35138 6880 36080 6886
rect 35138 6804 36030 6880
rect 35062 6798 36030 6804
rect 36066 6798 36080 6880
rect 45672 6886 46690 6894
rect 35062 6766 36080 6798
rect 37894 6806 38920 6834
rect 29968 6614 30910 6622
rect 29870 6584 30910 6614
rect 29870 5178 29992 6584
rect 33194 5178 33326 6684
rect 29476 5154 31312 5178
rect 29476 5120 29524 5154
rect 29892 5120 29982 5154
rect 30350 5120 30440 5154
rect 30808 5120 30898 5154
rect 31266 5120 31312 5154
rect 29476 5102 31312 5120
rect 31890 5161 33744 5178
rect 31890 5127 31951 5161
rect 32319 5127 32409 5161
rect 32777 5127 32867 5161
rect 33235 5127 33325 5161
rect 33693 5127 33744 5161
rect 29870 4970 29992 5102
rect 31890 5090 33744 5127
rect 29870 4914 29990 4970
rect 22666 4878 24664 4910
rect 28252 4888 29990 4914
rect 18551 4772 18568 4830
rect 22666 4780 24670 4878
rect 28252 4830 29084 4888
rect 29062 4822 29084 4830
rect 29150 4830 29990 4888
rect 33194 4910 33326 5090
rect 35062 4910 35192 6766
rect 37894 6720 37926 6806
rect 37966 6720 38842 6806
rect 38882 6720 38920 6806
rect 42906 6784 43942 6806
rect 42906 6778 43872 6784
rect 40408 6760 41438 6764
rect 37894 6702 38920 6720
rect 40398 6728 41438 6760
rect 40398 6720 41350 6728
rect 38784 4914 38916 6702
rect 40398 6614 40428 6720
rect 40496 6622 41350 6720
rect 41418 6622 41438 6728
rect 42906 6706 42962 6778
rect 42996 6706 43872 6778
rect 43908 6706 43942 6784
rect 42906 6684 43942 6706
rect 45672 6804 45712 6886
rect 45748 6880 46690 6886
rect 45748 6804 46640 6880
rect 45672 6798 46640 6804
rect 46676 6798 46690 6880
rect 56200 6886 57218 6894
rect 45672 6766 46690 6798
rect 48504 6806 49530 6834
rect 40496 6614 41438 6622
rect 40398 6584 41438 6614
rect 40398 5178 40520 6584
rect 43804 5178 43936 6684
rect 40004 5154 41840 5178
rect 40004 5120 40052 5154
rect 40420 5120 40510 5154
rect 40878 5120 40968 5154
rect 41336 5120 41426 5154
rect 41794 5120 41840 5154
rect 40004 5102 41840 5120
rect 42500 5161 44354 5178
rect 42500 5127 42561 5161
rect 42929 5127 43019 5161
rect 43387 5127 43477 5161
rect 43845 5127 43935 5161
rect 44303 5127 44354 5161
rect 40398 4970 40520 5102
rect 42500 5090 44354 5127
rect 40398 4914 40518 4970
rect 33194 4878 35192 4910
rect 38780 4886 40518 4914
rect 29150 4822 29176 4830
rect 18454 4142 18568 4772
rect 18454 4102 18472 4142
rect 18556 4102 18568 4142
rect 23566 4708 23784 4780
rect 23566 4548 23611 4708
rect 23748 4548 23784 4708
rect 21629 4122 21872 4136
rect 23566 4130 23784 4548
rect 18454 4088 18568 4102
rect 19550 4088 19618 4108
rect 11557 4044 12008 4078
rect 12042 4044 12060 4078
rect 11557 4033 12060 4044
rect 10854 4026 12060 4033
rect 12954 4034 13198 4050
rect 12954 3988 13018 4034
rect 13124 3988 13198 4034
rect 12954 3926 13198 3988
rect 12954 3880 13010 3926
rect 13116 3880 13198 3926
rect 12954 3770 13198 3880
rect 18446 4046 18582 4056
rect 18446 4006 18472 4046
rect 18552 4006 18582 4046
rect 18446 3940 18582 4006
rect 18446 3900 18474 3940
rect 18554 3900 18582 3940
rect 18446 3770 18582 3900
rect 19550 4054 19568 4088
rect 19602 4054 19618 4088
rect 12954 3590 18596 3770
rect 19550 3747 19618 4054
rect 21629 4103 22320 4122
rect 21629 4008 21653 4103
rect 21840 4096 22320 4103
rect 21840 4078 22668 4096
rect 23566 4094 23592 4130
rect 23732 4094 23784 4130
rect 23566 4080 23784 4094
rect 29062 4142 29176 4822
rect 33194 4780 35198 4878
rect 38780 4830 39612 4886
rect 39590 4796 39612 4830
rect 39688 4830 40518 4886
rect 43804 4910 43936 5090
rect 45672 4910 45802 6766
rect 48504 6720 48536 6806
rect 48576 6720 49452 6806
rect 49492 6720 49530 6806
rect 53434 6784 54470 6806
rect 53434 6778 54400 6784
rect 51018 6760 52048 6764
rect 48504 6702 49530 6720
rect 51008 6728 52048 6760
rect 51008 6720 51960 6728
rect 49394 4914 49526 6702
rect 51008 6614 51038 6720
rect 51106 6622 51960 6720
rect 52028 6622 52048 6728
rect 53434 6706 53490 6778
rect 53524 6706 54400 6778
rect 54436 6706 54470 6784
rect 53434 6684 54470 6706
rect 56200 6804 56240 6886
rect 56276 6880 57218 6886
rect 56276 6804 57168 6880
rect 56200 6798 57168 6804
rect 57204 6798 57218 6880
rect 56200 6766 57218 6798
rect 59032 6806 60058 6834
rect 51106 6614 52048 6622
rect 51008 6584 52048 6614
rect 51008 5178 51130 6584
rect 54332 5178 54464 6684
rect 50614 5154 52450 5178
rect 50614 5120 50662 5154
rect 51030 5120 51120 5154
rect 51488 5120 51578 5154
rect 51946 5120 52036 5154
rect 52404 5120 52450 5154
rect 50614 5102 52450 5120
rect 53028 5161 54882 5178
rect 53028 5127 53089 5161
rect 53457 5127 53547 5161
rect 53915 5127 54005 5161
rect 54373 5127 54463 5161
rect 54831 5127 54882 5161
rect 51008 4970 51130 5102
rect 53028 5090 54882 5127
rect 51008 4914 51128 4970
rect 43804 4878 45802 4910
rect 49390 4898 51128 4914
rect 39688 4796 39704 4830
rect 29062 4102 29080 4142
rect 29164 4102 29176 4142
rect 34094 4694 34312 4780
rect 34094 4532 34118 4694
rect 34290 4532 34312 4694
rect 34094 4130 34312 4532
rect 32108 4112 32799 4123
rect 29062 4088 29176 4102
rect 30158 4088 30227 4108
rect 21840 4044 22616 4078
rect 22650 4044 22668 4078
rect 21840 4026 22668 4044
rect 23562 4034 23806 4050
rect 21840 4008 22320 4026
rect 21629 3985 22320 4008
rect 23562 3988 23626 4034
rect 23732 3988 23806 4034
rect 23562 3926 23806 3988
rect 23562 3880 23618 3926
rect 23724 3880 23806 3926
rect 23562 3770 23806 3880
rect 29054 4046 29190 4056
rect 29054 4006 29080 4046
rect 29160 4006 29190 4046
rect 29054 3940 29190 4006
rect 29054 3900 29082 3940
rect 29162 3900 29190 3940
rect 29054 3770 29190 3900
rect 30158 4054 30176 4088
rect 30210 4054 30227 4088
rect 30158 3794 30227 4054
rect 32108 3997 32117 4112
rect 32324 4097 32799 4112
rect 32324 4096 33147 4097
rect 32324 4078 33196 4096
rect 34094 4094 34120 4130
rect 34260 4094 34312 4130
rect 34094 4080 34312 4094
rect 39590 4142 39704 4796
rect 43804 4780 45808 4878
rect 49390 4830 50212 4898
rect 50200 4826 50212 4830
rect 50300 4830 51128 4898
rect 54332 4910 54464 5090
rect 56200 4910 56330 6766
rect 59032 6720 59064 6806
rect 59104 6720 59980 6806
rect 60020 6720 60058 6806
rect 61546 6760 62576 6764
rect 59032 6702 60058 6720
rect 61536 6728 62576 6760
rect 61536 6720 62488 6728
rect 59922 4914 60054 6702
rect 61536 6614 61566 6720
rect 61634 6622 62488 6720
rect 62556 6622 62576 6728
rect 61634 6614 62576 6622
rect 61536 6584 62576 6614
rect 61536 5178 61658 6584
rect 61142 5154 62978 5178
rect 61142 5120 61190 5154
rect 61558 5120 61648 5154
rect 62016 5120 62106 5154
rect 62474 5120 62564 5154
rect 62932 5120 62978 5154
rect 61142 5102 62978 5120
rect 61536 4970 61658 5102
rect 61536 4914 61656 4970
rect 54332 4878 56330 4910
rect 59918 4896 61656 4914
rect 50300 4826 50314 4830
rect 44704 4740 44922 4780
rect 44704 4562 44746 4740
rect 44888 4562 44922 4740
rect 39590 4102 39608 4142
rect 39692 4102 39704 4142
rect 42782 4178 43384 4214
rect 39590 4088 39704 4102
rect 40686 4088 40754 4110
rect 32324 4044 33144 4078
rect 33178 4044 33196 4078
rect 32324 4027 33196 4044
rect 32324 3997 32799 4027
rect 33142 4026 33196 4027
rect 34090 4034 34334 4050
rect 32108 3986 32799 3997
rect 34090 3988 34154 4034
rect 34260 3988 34334 4034
rect 34090 3926 34334 3988
rect 34090 3880 34146 3926
rect 34252 3880 34334 3926
rect 19503 3662 19677 3747
rect 12954 3584 13198 3590
rect 16222 2976 16514 3590
rect 19503 3582 19533 3662
rect 19637 3582 19677 3662
rect 23562 3590 29204 3770
rect 30004 3696 30385 3794
rect 23562 3584 23806 3590
rect 19503 3544 19677 3582
rect 26830 2976 27122 3590
rect 30004 3558 30133 3696
rect 30272 3558 30385 3696
rect 34090 3770 34334 3880
rect 39582 4046 39718 4056
rect 39582 4006 39608 4046
rect 39688 4006 39718 4046
rect 39582 3940 39718 4006
rect 39582 3900 39610 3940
rect 39690 3900 39718 3940
rect 39582 3770 39718 3900
rect 40686 4054 40704 4088
rect 40738 4054 40754 4088
rect 34090 3590 39732 3770
rect 40686 3750 40754 4054
rect 42782 3854 42806 4178
rect 42960 4096 43384 4178
rect 44704 4130 44922 4562
rect 42960 4078 43806 4096
rect 44704 4094 44730 4130
rect 44870 4094 44922 4130
rect 44704 4080 44922 4094
rect 50200 4142 50314 4826
rect 54332 4780 56336 4878
rect 59918 4830 60745 4896
rect 60728 4804 60745 4830
rect 60821 4830 61656 4896
rect 60821 4804 60842 4830
rect 55232 4612 55450 4780
rect 55232 4392 55246 4612
rect 55425 4392 55450 4612
rect 50200 4102 50218 4142
rect 50302 4102 50314 4142
rect 53268 4184 53844 4238
rect 50200 4088 50314 4102
rect 51296 4088 51364 4108
rect 42960 4044 43754 4078
rect 43788 4044 43806 4078
rect 42960 4026 43806 4044
rect 44700 4034 44944 4050
rect 42960 3854 43384 4026
rect 42782 3830 43384 3854
rect 44700 3988 44764 4034
rect 44870 3988 44944 4034
rect 44700 3926 44944 3988
rect 44700 3880 44756 3926
rect 44862 3880 44944 3926
rect 44700 3770 44944 3880
rect 50192 4046 50328 4056
rect 50192 4006 50218 4046
rect 50298 4006 50328 4046
rect 50192 3940 50328 4006
rect 50192 3900 50220 3940
rect 50300 3900 50328 3940
rect 50192 3770 50328 3900
rect 51296 4054 51314 4088
rect 51348 4054 51364 4088
rect 51296 3782 51364 4054
rect 53268 3910 53318 4184
rect 53780 4096 53844 4184
rect 55232 4130 55450 4392
rect 53780 4078 54334 4096
rect 55232 4094 55258 4130
rect 55398 4094 55450 4130
rect 55232 4080 55450 4094
rect 60728 4142 60842 4804
rect 60728 4102 60746 4142
rect 60830 4102 60842 4142
rect 60728 4088 60842 4102
rect 61824 4088 61894 4108
rect 53780 4044 54282 4078
rect 54316 4044 54334 4078
rect 53780 4026 54334 4044
rect 55228 4034 55472 4050
rect 53780 3910 53844 4026
rect 53268 3860 53844 3910
rect 55228 3988 55292 4034
rect 55398 3988 55472 4034
rect 55228 3926 55472 3988
rect 55228 3880 55284 3926
rect 55390 3880 55472 3926
rect 40564 3642 40956 3750
rect 34090 3584 34334 3590
rect 30004 3454 30385 3558
rect 30158 3453 30227 3454
rect 37358 2976 37650 3590
rect 40564 3478 40672 3642
rect 40838 3478 40956 3642
rect 44700 3590 50342 3770
rect 51178 3722 51504 3782
rect 44700 3584 44944 3590
rect 40564 3368 40956 3478
rect 47968 2976 48260 3590
rect 51178 3460 51212 3722
rect 51468 3460 51504 3722
rect 55228 3770 55472 3880
rect 60720 4046 60856 4056
rect 60720 4006 60746 4046
rect 60826 4006 60856 4046
rect 60720 3940 60856 4006
rect 60720 3900 60748 3940
rect 60828 3900 60856 3940
rect 60720 3770 60856 3900
rect 61824 4054 61842 4088
rect 61876 4054 61894 4088
rect 61824 3790 61894 4054
rect 55228 3590 60870 3770
rect 61730 3752 62004 3790
rect 55228 3584 55472 3590
rect 51178 3426 51504 3460
rect 58496 2976 58788 3590
rect 61730 3586 61786 3752
rect 61960 3586 62004 3752
rect 61730 3298 62004 3586
rect 14366 2970 19074 2976
rect 14366 2962 17164 2970
rect 14366 2958 16256 2962
rect 14366 2862 14422 2958
rect 14470 2950 16256 2958
rect 14470 2862 15338 2950
rect 14366 2854 15338 2862
rect 15386 2866 16256 2950
rect 16304 2874 17164 2962
rect 17212 2964 19074 2970
rect 17212 2874 18070 2964
rect 16304 2868 18070 2874
rect 18118 2868 19002 2964
rect 19050 2868 19074 2964
rect 16304 2866 19074 2868
rect 15386 2854 19074 2866
rect 14366 2844 19074 2854
rect 24974 2970 29682 2976
rect 24974 2962 27772 2970
rect 24974 2958 26864 2962
rect 24974 2862 25030 2958
rect 25078 2950 26864 2958
rect 25078 2862 25946 2950
rect 24974 2854 25946 2862
rect 25994 2866 26864 2950
rect 26912 2874 27772 2962
rect 27820 2964 29682 2970
rect 27820 2874 28678 2964
rect 26912 2868 28678 2874
rect 28726 2868 29610 2964
rect 29658 2868 29682 2964
rect 26912 2866 29682 2868
rect 25994 2854 29682 2866
rect 24974 2844 29682 2854
rect 35502 2970 40210 2976
rect 35502 2962 38300 2970
rect 35502 2958 37392 2962
rect 35502 2862 35558 2958
rect 35606 2950 37392 2958
rect 35606 2862 36474 2950
rect 35502 2854 36474 2862
rect 36522 2866 37392 2950
rect 37440 2874 38300 2962
rect 38348 2964 40210 2970
rect 38348 2874 39206 2964
rect 37440 2868 39206 2874
rect 39254 2868 40138 2964
rect 40186 2868 40210 2964
rect 37440 2866 40210 2868
rect 36522 2854 40210 2866
rect 35502 2844 40210 2854
rect 46112 2970 50820 2976
rect 46112 2962 48910 2970
rect 46112 2958 48002 2962
rect 46112 2862 46168 2958
rect 46216 2950 48002 2958
rect 46216 2862 47084 2950
rect 46112 2854 47084 2862
rect 47132 2866 48002 2950
rect 48050 2874 48910 2962
rect 48958 2964 50820 2970
rect 48958 2874 49816 2964
rect 48050 2868 49816 2874
rect 49864 2868 50748 2964
rect 50796 2868 50820 2964
rect 48050 2866 50820 2868
rect 47132 2854 50820 2866
rect 46112 2844 50820 2854
rect 56640 2970 61348 2976
rect 56640 2962 59438 2970
rect 56640 2958 58530 2962
rect 56640 2862 56696 2958
rect 56744 2950 58530 2958
rect 56744 2862 57612 2950
rect 56640 2854 57612 2862
rect 57660 2866 58530 2950
rect 58578 2874 59438 2962
rect 59486 2964 61348 2970
rect 59486 2874 60344 2964
rect 58578 2868 60344 2874
rect 60392 2868 61276 2964
rect 61324 2868 61348 2964
rect 58578 2866 61348 2868
rect 57660 2854 61348 2866
rect 56640 2844 61348 2854
rect 16222 2834 16514 2844
rect 26830 2834 27122 2844
rect 37358 2834 37650 2844
rect 47968 2834 48260 2844
rect 58496 2834 58788 2844
rect 14802 2786 19556 2792
rect 14802 2780 19440 2786
rect 14802 2768 16696 2780
rect 14802 2756 15778 2768
rect 14802 2646 14854 2756
rect 14924 2658 15778 2756
rect 15848 2758 16696 2768
rect 16766 2758 17620 2780
rect 15848 2658 16684 2758
rect 16798 2670 17620 2758
rect 17690 2768 19440 2780
rect 17690 2670 18544 2768
rect 14924 2650 16684 2658
rect 16798 2658 18544 2670
rect 18614 2676 19440 2768
rect 19510 2676 19556 2786
rect 18614 2658 19556 2676
rect 16798 2650 19556 2658
rect 14924 2646 19556 2650
rect 14802 2628 19556 2646
rect 25410 2786 30164 2792
rect 25410 2780 30048 2786
rect 25410 2768 27304 2780
rect 25410 2756 26386 2768
rect 25410 2646 25462 2756
rect 25532 2658 26386 2756
rect 26456 2758 27304 2768
rect 27374 2758 28228 2780
rect 26456 2658 27292 2758
rect 27406 2670 28228 2758
rect 28298 2768 30048 2780
rect 28298 2670 29152 2768
rect 25532 2650 27292 2658
rect 27406 2658 29152 2670
rect 29222 2676 30048 2768
rect 30118 2676 30164 2786
rect 29222 2658 30164 2676
rect 27406 2650 30164 2658
rect 25532 2646 30164 2650
rect 25410 2628 30164 2646
rect 35938 2786 40692 2792
rect 35938 2780 40576 2786
rect 35938 2768 37832 2780
rect 35938 2756 36914 2768
rect 35938 2646 35990 2756
rect 36060 2658 36914 2756
rect 36984 2758 37832 2768
rect 37902 2758 38756 2780
rect 36984 2658 37820 2758
rect 37934 2670 38756 2758
rect 38826 2768 40576 2780
rect 38826 2670 39680 2768
rect 36060 2650 37820 2658
rect 37934 2658 39680 2670
rect 39750 2676 40576 2768
rect 40646 2676 40692 2786
rect 39750 2658 40692 2676
rect 37934 2650 40692 2658
rect 36060 2646 40692 2650
rect 35938 2628 40692 2646
rect 46548 2786 51302 2792
rect 46548 2780 51186 2786
rect 46548 2768 48442 2780
rect 46548 2756 47524 2768
rect 46548 2646 46600 2756
rect 46670 2658 47524 2756
rect 47594 2758 48442 2768
rect 48512 2758 49366 2780
rect 47594 2658 48430 2758
rect 48544 2670 49366 2758
rect 49436 2768 51186 2780
rect 49436 2670 50290 2768
rect 46670 2650 48430 2658
rect 48544 2658 50290 2670
rect 50360 2676 51186 2768
rect 51256 2676 51302 2786
rect 50360 2658 51302 2676
rect 48544 2650 51302 2658
rect 46670 2646 51302 2650
rect 46548 2628 51302 2646
rect 57076 2786 61830 2792
rect 57076 2780 61714 2786
rect 57076 2768 58970 2780
rect 57076 2756 58052 2768
rect 57076 2646 57128 2756
rect 57198 2658 58052 2756
rect 58122 2758 58970 2768
rect 59040 2758 59894 2780
rect 58122 2658 58958 2758
rect 59072 2670 59894 2758
rect 59964 2768 61714 2780
rect 59964 2670 60818 2768
rect 57198 2650 58958 2658
rect 59072 2658 60818 2670
rect 60888 2676 61714 2768
rect 61784 2676 61830 2786
rect 60888 2658 61830 2676
rect 59072 2650 61830 2658
rect 57198 2646 61830 2650
rect 57076 2628 61830 2646
rect 12867 615 61802 648
rect 12867 581 14491 615
rect 14859 581 14949 615
rect 15317 581 15407 615
rect 15775 581 15865 615
rect 16233 581 16323 615
rect 16691 581 16781 615
rect 17149 581 17239 615
rect 17607 581 17697 615
rect 18065 581 18155 615
rect 18523 581 18613 615
rect 18981 581 19071 615
rect 19439 581 25099 615
rect 25467 581 25557 615
rect 25925 581 26015 615
rect 26383 581 26473 615
rect 26841 581 26931 615
rect 27299 581 27389 615
rect 27757 581 27847 615
rect 28215 581 28305 615
rect 28673 581 28763 615
rect 29131 581 29221 615
rect 29589 581 29679 615
rect 30047 581 35627 615
rect 35995 581 36085 615
rect 36453 581 36543 615
rect 36911 581 37001 615
rect 37369 581 37459 615
rect 37827 581 37917 615
rect 38285 581 38375 615
rect 38743 581 38833 615
rect 39201 581 39291 615
rect 39659 581 39749 615
rect 40117 581 40207 615
rect 40575 581 46237 615
rect 46605 581 46695 615
rect 47063 581 47153 615
rect 47521 581 47611 615
rect 47979 581 48069 615
rect 48437 581 48527 615
rect 48895 581 48985 615
rect 49353 581 49443 615
rect 49811 581 49901 615
rect 50269 581 50359 615
rect 50727 581 50817 615
rect 51185 581 56765 615
rect 57133 581 57223 615
rect 57591 581 57681 615
rect 58049 581 58139 615
rect 58507 581 58597 615
rect 58965 581 59055 615
rect 59423 581 59513 615
rect 59881 581 59971 615
rect 60339 581 60429 615
rect 60797 581 60887 615
rect 61255 581 61345 615
rect 61713 581 61802 615
rect 12867 566 61802 581
rect 12867 562 14546 566
rect 24592 562 25154 566
rect 35120 562 35682 566
rect 45730 562 46292 566
rect 56258 562 56820 566
rect 18322 504 18498 532
rect 18322 470 18344 504
rect 18446 470 18498 504
rect 18322 362 18498 470
rect 28930 504 29106 532
rect 28930 470 28952 504
rect 29054 470 29106 504
rect 28930 362 29106 470
rect 39458 504 39634 532
rect 39458 470 39480 504
rect 39582 470 39634 504
rect 39458 362 39634 470
rect 50068 504 50244 532
rect 50068 470 50090 504
rect 50192 470 50244 504
rect 50068 362 50244 470
rect 60596 504 60772 532
rect 60596 470 60618 504
rect 60720 470 60772 504
rect 60596 362 60772 470
rect 10548 278 63264 362
rect 10548 272 17148 278
rect 10548 164 14372 272
rect 14486 256 16208 272
rect 14486 164 15318 256
rect 10548 148 15318 164
rect 15432 164 16208 256
rect 16322 254 17148 272
rect 16322 164 16684 254
rect 15432 148 16684 164
rect 10548 146 16684 148
rect 16798 170 17148 254
rect 17262 272 18970 278
rect 17262 170 18076 272
rect 16798 164 18076 170
rect 18190 170 18970 272
rect 19084 272 27756 278
rect 19084 170 24980 272
rect 18190 164 24980 170
rect 25094 256 26816 272
rect 25094 164 25926 256
rect 16798 148 25926 164
rect 26040 164 26816 256
rect 26930 254 27756 272
rect 26930 164 27292 254
rect 26040 148 27292 164
rect 16798 146 27292 148
rect 27406 170 27756 254
rect 27870 272 29578 278
rect 27870 170 28684 272
rect 27406 164 28684 170
rect 28798 170 29578 272
rect 29692 272 38284 278
rect 29692 170 35508 272
rect 28798 164 35508 170
rect 35622 256 37344 272
rect 35622 164 36454 256
rect 27406 148 36454 164
rect 36568 164 37344 256
rect 37458 254 38284 272
rect 37458 164 37820 254
rect 36568 148 37820 164
rect 27406 146 37820 148
rect 37934 170 38284 254
rect 38398 272 40106 278
rect 38398 170 39212 272
rect 37934 164 39212 170
rect 39326 170 40106 272
rect 40220 272 48894 278
rect 40220 170 46118 272
rect 39326 164 46118 170
rect 46232 256 47954 272
rect 46232 164 47064 256
rect 37934 148 47064 164
rect 47178 164 47954 256
rect 48068 254 48894 272
rect 48068 164 48430 254
rect 47178 148 48430 164
rect 37934 146 48430 148
rect 48544 170 48894 254
rect 49008 272 50716 278
rect 49008 170 49822 272
rect 48544 164 49822 170
rect 49936 170 50716 272
rect 50830 272 59422 278
rect 50830 170 56646 272
rect 49936 164 56646 170
rect 56760 256 58482 272
rect 56760 164 57592 256
rect 48544 148 57592 164
rect 57706 164 58482 256
rect 58596 254 59422 272
rect 58596 164 58958 254
rect 57706 148 58958 164
rect 48544 146 58958 148
rect 59072 170 59422 254
rect 59536 272 61244 278
rect 59536 170 60350 272
rect 59072 164 60350 170
rect 60464 170 61244 272
rect 61358 170 63264 278
rect 60464 164 63264 170
rect 59072 146 63264 164
rect 10548 -128 63264 146
<< via1 >>
rect 16320 7686 16374 7696
rect 13496 7580 13608 7670
rect 16320 7606 16374 7686
rect 26928 7686 26982 7696
rect 24104 7580 24216 7670
rect 26928 7606 26982 7686
rect 37456 7686 37510 7696
rect 34632 7580 34744 7670
rect 37456 7606 37510 7686
rect 48066 7686 48120 7696
rect 45242 7580 45354 7670
rect 48066 7606 48120 7686
rect 58594 7686 58648 7696
rect 55770 7580 55882 7670
rect 58594 7606 58648 7686
rect 15765 7185 15972 7304
rect 13500 7022 13508 7094
rect 13508 7022 13544 7094
rect 13544 7022 13606 7094
rect 13500 7002 13606 7022
rect 16318 7006 16328 7088
rect 16328 7006 16372 7088
rect 16318 6998 16372 7006
rect 26375 7180 26582 7299
rect 24108 7022 24116 7094
rect 24116 7022 24152 7094
rect 24152 7022 24214 7094
rect 24108 7002 24214 7022
rect 26926 7006 26936 7088
rect 26936 7006 26980 7088
rect 26926 6998 26980 7006
rect 36904 7180 37111 7299
rect 34636 7022 34644 7094
rect 34644 7022 34680 7094
rect 34680 7022 34742 7094
rect 34636 7002 34742 7022
rect 37454 7006 37464 7088
rect 37464 7006 37508 7088
rect 37454 6998 37508 7006
rect 47487 7180 47694 7299
rect 45246 7022 45254 7094
rect 45254 7022 45290 7094
rect 45290 7022 45352 7094
rect 45246 7002 45352 7022
rect 48064 7006 48074 7088
rect 48074 7006 48118 7088
rect 48064 6998 48118 7006
rect 58057 7194 58264 7313
rect 55774 7022 55782 7094
rect 55782 7022 55818 7094
rect 55818 7022 55880 7094
rect 55774 7002 55880 7022
rect 58592 7006 58602 7088
rect 58602 7006 58646 7088
rect 58592 6998 58646 7006
rect 12996 4499 13134 4636
rect 10871 4033 11557 4090
rect 18476 4772 18551 4869
rect 29084 4822 29150 4888
rect 23611 4548 23748 4708
rect 21653 4008 21840 4103
rect 39612 4796 39688 4886
rect 34118 4532 34290 4694
rect 32117 3997 32324 4112
rect 50212 4826 50300 4898
rect 44746 4562 44888 4740
rect 19533 3582 19637 3662
rect 30133 3558 30272 3696
rect 42806 3854 42960 4178
rect 60745 4804 60821 4896
rect 55246 4392 55425 4612
rect 53318 3910 53780 4184
rect 40672 3478 40838 3642
rect 51212 3460 51468 3722
rect 61786 3586 61960 3752
rect 16684 2670 16696 2758
rect 16696 2670 16766 2758
rect 16766 2670 16798 2758
rect 16684 2650 16798 2670
rect 27292 2670 27304 2758
rect 27304 2670 27374 2758
rect 27374 2670 27406 2758
rect 27292 2650 27406 2670
rect 37820 2670 37832 2758
rect 37832 2670 37902 2758
rect 37902 2670 37934 2758
rect 37820 2650 37934 2670
rect 48430 2670 48442 2758
rect 48442 2670 48512 2758
rect 48512 2670 48544 2758
rect 48430 2650 48544 2670
rect 58958 2670 58970 2758
rect 58970 2670 59040 2758
rect 59040 2670 59072 2758
rect 58958 2650 59072 2670
rect 16684 146 16798 254
rect 27292 146 27406 254
rect 37820 146 37934 254
rect 48430 146 48544 254
rect 58958 146 59072 254
<< metal2 >>
rect 4840 14270 10391 14273
rect 64015 14270 65864 14307
rect 4840 14124 65864 14270
rect 4840 13083 64676 14124
rect 65695 13083 65864 14124
rect 4840 12949 65864 13083
rect 4840 12942 64321 12949
rect 4840 3694 6567 12942
rect 10168 11148 64271 11154
rect 8738 9826 64271 11148
rect 8738 4282 10278 9826
rect 13474 7670 13646 7764
rect 13474 7580 13496 7670
rect 13608 7580 13646 7670
rect 13474 7094 13646 7580
rect 16304 7696 16390 7772
rect 16304 7606 16320 7696
rect 16374 7606 16390 7696
rect 15722 7332 16011 7351
rect 15722 7161 15741 7332
rect 15994 7161 16011 7332
rect 15722 7142 16011 7161
rect 13474 7002 13500 7094
rect 13606 7002 13646 7094
rect 13474 6962 13646 7002
rect 16304 7088 16390 7606
rect 16304 6998 16318 7088
rect 16372 6998 16390 7088
rect 16304 6966 16390 6998
rect 24082 7670 24254 7764
rect 24082 7580 24104 7670
rect 24216 7580 24254 7670
rect 24082 7094 24254 7580
rect 26912 7696 26998 7772
rect 26912 7606 26928 7696
rect 26982 7606 26998 7696
rect 26332 7327 26621 7346
rect 26332 7156 26351 7327
rect 26604 7156 26621 7327
rect 26332 7137 26621 7156
rect 24082 7002 24108 7094
rect 24214 7002 24254 7094
rect 24082 6962 24254 7002
rect 26912 7088 26998 7606
rect 26912 6998 26926 7088
rect 26980 6998 26998 7088
rect 26912 6966 26998 6998
rect 34610 7670 34782 7764
rect 34610 7580 34632 7670
rect 34744 7580 34782 7670
rect 34610 7094 34782 7580
rect 37440 7696 37526 7772
rect 37440 7606 37456 7696
rect 37510 7606 37526 7696
rect 36861 7327 37150 7346
rect 36861 7156 36880 7327
rect 37133 7156 37150 7327
rect 36861 7137 37150 7156
rect 34610 7002 34636 7094
rect 34742 7002 34782 7094
rect 34610 6962 34782 7002
rect 37440 7088 37526 7606
rect 37440 6998 37454 7088
rect 37508 6998 37526 7088
rect 37440 6966 37526 6998
rect 45220 7670 45392 7764
rect 45220 7580 45242 7670
rect 45354 7580 45392 7670
rect 45220 7094 45392 7580
rect 48050 7696 48136 7772
rect 48050 7606 48066 7696
rect 48120 7606 48136 7696
rect 47444 7327 47733 7346
rect 47444 7156 47463 7327
rect 47716 7156 47733 7327
rect 47444 7137 47733 7156
rect 45220 7002 45246 7094
rect 45352 7002 45392 7094
rect 45220 6962 45392 7002
rect 48050 7088 48136 7606
rect 48050 6998 48064 7088
rect 48118 6998 48136 7088
rect 48050 6966 48136 6998
rect 55748 7670 55920 7764
rect 55748 7580 55770 7670
rect 55882 7580 55920 7670
rect 55748 7094 55920 7580
rect 58578 7696 58664 7772
rect 58578 7606 58594 7696
rect 58648 7606 58664 7696
rect 58014 7341 58303 7360
rect 58014 7170 58033 7341
rect 58286 7170 58303 7341
rect 58014 7151 58303 7170
rect 55748 7002 55774 7094
rect 55880 7002 55920 7094
rect 55748 6962 55920 7002
rect 58578 7088 58664 7606
rect 58578 6998 58592 7088
rect 58646 6998 58664 7088
rect 58578 6966 58664 6998
rect 18450 4884 18573 4911
rect 18450 4768 18469 4884
rect 18554 4768 18573 4884
rect 29058 4910 29182 4924
rect 29058 4812 29076 4910
rect 29166 4812 29182 4910
rect 29058 4796 29182 4812
rect 39570 4898 39724 4920
rect 39570 4802 39594 4898
rect 39700 4802 39724 4898
rect 50198 4908 50320 4920
rect 50198 4824 50210 4908
rect 50306 4824 50320 4908
rect 50198 4812 50320 4824
rect 60717 4901 60864 4930
rect 39570 4796 39612 4802
rect 39688 4796 39724 4802
rect 39570 4776 39724 4796
rect 60717 4796 60739 4901
rect 60848 4796 60864 4901
rect 60717 4775 60864 4796
rect 18450 4751 18573 4768
rect 44668 4740 53564 4772
rect 32043 4725 32367 4730
rect 23526 4708 32367 4725
rect 12913 4636 21875 4662
rect 12913 4499 12996 4636
rect 13134 4499 21875 4636
rect 23526 4548 23611 4708
rect 23748 4548 32367 4708
rect 23526 4504 32367 4548
rect 12913 4451 21875 4499
rect 8738 4194 11020 4282
rect 8738 4090 12065 4194
rect 8738 4033 10871 4090
rect 11557 4033 12065 4090
rect 8738 3930 12065 4033
rect 21629 4103 21875 4451
rect 21629 4008 21653 4103
rect 21840 4008 21875 4103
rect 21629 3985 21875 4008
rect 32043 4112 32367 4504
rect 34066 4694 42996 4724
rect 34066 4532 34118 4694
rect 34290 4532 42996 4694
rect 34066 4500 42996 4532
rect 44668 4562 44746 4740
rect 44888 4562 53564 4740
rect 63686 4674 64271 9826
rect 44668 4510 53564 4562
rect 55170 4612 64271 4674
rect 32043 3997 32117 4112
rect 32324 3997 32367 4112
rect 8738 3924 11020 3930
rect 32043 3804 32367 3997
rect 42780 4178 42992 4500
rect 42780 3854 42806 4178
rect 42960 3854 42992 4178
rect 53268 4238 53560 4510
rect 55170 4392 55246 4612
rect 55425 4392 64271 4612
rect 55170 4302 64271 4392
rect 63686 4299 64271 4302
rect 53268 4184 53844 4238
rect 53268 3910 53318 4184
rect 53780 3910 53844 4184
rect 53268 3860 53844 3910
rect 42780 3834 42992 3854
rect 30004 3696 30385 3794
rect 4840 3688 8961 3694
rect 4840 3662 19677 3688
rect 4840 3582 19533 3662
rect 19637 3582 19677 3662
rect 4840 3427 19677 3582
rect 30004 3681 30133 3696
rect 30272 3681 30385 3696
rect 30004 3471 30025 3681
rect 30360 3471 30385 3681
rect 30004 3454 30385 3471
rect 40564 3642 40956 3750
rect 40564 3506 40672 3642
rect 40838 3506 40956 3642
rect 4840 3232 8961 3427
rect 40564 3396 40600 3506
rect 40914 3396 40956 3506
rect 51178 3722 51504 3782
rect 51178 3460 51212 3722
rect 51468 3644 51504 3722
rect 51474 3478 51504 3644
rect 51468 3460 51504 3478
rect 51178 3426 51504 3460
rect 61730 3752 62004 3790
rect 61730 3586 61786 3752
rect 61960 3586 62004 3752
rect 61730 3514 62004 3586
rect 40564 3368 40956 3396
rect 61730 3310 61748 3514
rect 61914 3310 62004 3514
rect 61730 3298 62004 3310
rect 4840 3209 6567 3232
rect 16662 2758 16844 2780
rect 16662 2650 16684 2758
rect 16798 2650 16844 2758
rect 16662 254 16844 2650
rect 16662 146 16684 254
rect 16798 146 16844 254
rect 16662 138 16844 146
rect 27270 2758 27452 2780
rect 27270 2650 27292 2758
rect 27406 2650 27452 2758
rect 27270 254 27452 2650
rect 27270 146 27292 254
rect 27406 146 27452 254
rect 27270 138 27452 146
rect 37798 2758 37980 2780
rect 37798 2650 37820 2758
rect 37934 2650 37980 2758
rect 37798 254 37980 2650
rect 37798 146 37820 254
rect 37934 146 37980 254
rect 37798 138 37980 146
rect 48408 2758 48590 2780
rect 48408 2650 48430 2758
rect 48544 2650 48590 2758
rect 48408 254 48590 2650
rect 48408 146 48430 254
rect 48544 146 48590 254
rect 48408 138 48590 146
rect 58936 2758 59118 2780
rect 58936 2650 58958 2758
rect 59072 2650 59118 2758
rect 58936 254 59118 2650
rect 58936 146 58958 254
rect 59072 146 59118 254
rect 58936 138 59118 146
<< via2 >>
rect 64676 13083 65695 14124
rect 15741 7304 15994 7332
rect 15741 7185 15765 7304
rect 15765 7185 15972 7304
rect 15972 7185 15994 7304
rect 15741 7161 15994 7185
rect 26351 7299 26604 7327
rect 26351 7180 26375 7299
rect 26375 7180 26582 7299
rect 26582 7180 26604 7299
rect 26351 7156 26604 7180
rect 36880 7299 37133 7327
rect 36880 7180 36904 7299
rect 36904 7180 37111 7299
rect 37111 7180 37133 7299
rect 36880 7156 37133 7180
rect 47463 7299 47716 7327
rect 47463 7180 47487 7299
rect 47487 7180 47694 7299
rect 47694 7180 47716 7299
rect 47463 7156 47716 7180
rect 58033 7313 58286 7341
rect 58033 7194 58057 7313
rect 58057 7194 58264 7313
rect 58264 7194 58286 7313
rect 58033 7170 58286 7194
rect 18469 4869 18554 4884
rect 18469 4772 18476 4869
rect 18476 4772 18551 4869
rect 18551 4772 18554 4869
rect 18469 4768 18554 4772
rect 29076 4888 29166 4910
rect 29076 4822 29084 4888
rect 29084 4822 29150 4888
rect 29150 4822 29166 4888
rect 29076 4812 29166 4822
rect 39594 4886 39700 4898
rect 39594 4802 39612 4886
rect 39612 4802 39688 4886
rect 39688 4802 39700 4886
rect 50210 4898 50306 4908
rect 50210 4826 50212 4898
rect 50212 4826 50300 4898
rect 50300 4826 50306 4898
rect 50210 4824 50306 4826
rect 60739 4896 60848 4901
rect 60739 4804 60745 4896
rect 60745 4804 60821 4896
rect 60821 4804 60848 4896
rect 60739 4796 60848 4804
rect 30025 3558 30133 3681
rect 30133 3558 30272 3681
rect 30272 3558 30360 3681
rect 30025 3471 30360 3558
rect 40600 3478 40672 3506
rect 40672 3478 40838 3506
rect 40838 3478 40914 3506
rect 40600 3396 40914 3478
rect 51216 3478 51468 3644
rect 51468 3478 51474 3644
rect 61748 3310 61914 3514
<< metal3 >>
rect 64563 14124 65878 14314
rect 64563 13083 64676 14124
rect 65695 13083 65878 14124
rect 15223 8687 58317 8750
rect 15223 8364 15282 8687
rect 15754 8364 58317 8687
rect 15223 8307 58317 8364
rect 15710 7332 16025 8307
rect 15710 7161 15741 7332
rect 15994 7161 16025 7332
rect 15710 7127 16025 7161
rect 26320 7327 26635 8307
rect 36848 7362 37163 8307
rect 36848 7331 37164 7362
rect 26320 7156 26351 7327
rect 26604 7156 26635 7327
rect 26320 7122 26635 7156
rect 36849 7327 37164 7331
rect 36849 7156 36880 7327
rect 37133 7156 37164 7327
rect 36849 7122 37164 7156
rect 47432 7327 47747 8307
rect 47432 7156 47463 7327
rect 47716 7156 47747 7327
rect 47432 7122 47747 7156
rect 58002 7341 58317 8307
rect 58002 7170 58033 7341
rect 58286 7170 58317 7341
rect 58002 7136 58317 7170
rect 64563 4943 65878 13083
rect 18440 4884 20927 4916
rect 18440 4768 18469 4884
rect 18554 4768 20927 4884
rect 29006 4910 31678 4936
rect 29006 4812 29076 4910
rect 29166 4812 31678 4910
rect 29006 4776 31678 4812
rect 39532 4898 42334 4936
rect 39532 4802 39594 4898
rect 39700 4802 42334 4898
rect 18440 4746 20927 4768
rect 20754 4150 20927 4746
rect 20708 3708 21009 4150
rect 20708 3681 30384 3708
rect 20708 3471 30025 3681
rect 30360 3471 30384 3681
rect 20708 3454 30384 3471
rect 31368 3544 31676 4776
rect 39532 4760 42334 4802
rect 50186 4908 53056 4938
rect 50186 4824 50210 4908
rect 50306 4824 53056 4908
rect 50186 4800 53056 4824
rect 60692 4901 65878 4943
rect 42060 3674 42332 4760
rect 42060 3644 51490 3674
rect 31368 3506 40950 3544
rect 20708 3448 21009 3454
rect 31368 3396 40600 3506
rect 40914 3396 40950 3506
rect 31368 3368 40950 3396
rect 42060 3478 51216 3644
rect 51474 3478 51490 3644
rect 52828 3540 53054 4800
rect 60692 4796 60739 4901
rect 60848 4796 65878 4901
rect 60692 4757 65878 4796
rect 64563 4687 65878 4757
rect 42060 3436 51490 3478
rect 52820 3514 61930 3540
rect 42060 3142 42332 3436
rect 52820 3310 61748 3514
rect 61914 3310 61930 3514
rect 52820 3292 61930 3310
rect 52828 3070 53054 3292
<< via3 >>
rect 15282 8364 15754 8687
<< metal4 >>
rect 15219 8710 15853 8773
rect 15219 8687 15292 8710
rect 15219 8364 15282 8687
rect 15219 8351 15292 8364
rect 15803 8351 15853 8710
rect 15219 8291 15853 8351
<< via4 >>
rect 15292 8687 15803 8710
rect 15292 8364 15754 8687
rect 15754 8364 15803 8687
rect 15292 8351 15803 8364
<< metal5 >>
rect 15038 8710 15935 8901
rect 15038 8351 15292 8710
rect 15803 8351 15935 8710
rect 15038 8238 15935 8351
<< labels >>
rlabel metal1 11774 7522 11994 7750 1 Vdd
port 1 n
rlabel metal1 15850 7238 15980 7288 1 Vctrl
port 3 n
rlabel metal1 14002 574 14094 644 1 vbn
port 8 n
rlabel metal1 16458 130 16616 246 1 Gnd
port 9 n
rlabel metal1 32910 7522 33130 7750 1 Vdd
port 1 n
rlabel metal1 36986 7238 37116 7288 1 Vctrl
port 3 n
rlabel metal1 35138 574 35230 644 1 vbn
port 8 n
rlabel metal1 37594 130 37752 246 1 Gnd
port 9 n
rlabel metal1 22382 7522 22602 7750 1 Vdd
port 1 n
rlabel metal1 26458 7238 26588 7288 1 Vctrl
port 3 n
rlabel metal1 24610 574 24702 644 1 vbn
port 8 n
rlabel metal1 27066 130 27224 246 1 Gnd
port 9 n
rlabel metal1 54048 7522 54268 7750 1 Vdd
port 1 n
rlabel via1 58124 7238 58254 7288 1 Vctrl
port 3 n
rlabel metal1 56276 574 56368 644 1 vbn
port 8 n
rlabel metal1 58732 130 58890 246 1 Gnd
port 9 n
rlabel metal1 43520 7522 43740 7750 1 Vdd
port 1 n
rlabel metal1 47596 7238 47726 7288 1 Vctrl
port 3 n
rlabel metal1 45748 574 45840 644 1 vbn
port 8 n
rlabel metal1 48204 130 48362 246 1 Gnd
port 9 n
rlabel metal1 58166 7252 58296 7302 1 Vctrl
port 3 n
rlabel metal2 8970 4110 10102 4746 1 inp
port 10 n
rlabel metal2 5148 4118 6280 4754 1 inn
port 11 n
<< end >>
