magic
tech sky130A
magscale 1 2
timestamp 1606531739
<< pwell >>
rect 168611 -27625 168750 -27565
<< locali >>
rect 165785 -25054 166173 -24622
rect 166421 -25054 166809 -24622
rect 167057 -25054 167445 -24622
rect 167693 -25054 168081 -24622
rect 168329 -25054 168717 -24622
rect 164438 -26674 165689 -25938
rect 146718 -27412 156544 -27258
rect 146718 -28390 156580 -27412
rect 166103 -27486 166491 -27054
rect 166739 -27486 167127 -27054
rect 167375 -27486 167763 -27054
rect 168011 -27486 168399 -27054
rect 165655 -28392 166532 -27614
rect 146718 -30726 146820 -30698
rect 156480 -30726 156580 -30698
rect 146718 -30732 156580 -30726
<< viali >>
rect 160358 -26118 164326 -26084
rect 160358 -26528 164326 -26494
rect 165785 -27486 165855 -27054
rect 168647 -27486 168717 -27054
rect 146820 -30726 156480 -30684
rect 157854 -30726 167514 -30684
<< metal1 >>
rect 156671 -25046 156781 -25001
rect 156671 -27139 156691 -25046
rect 156752 -27179 156781 -25046
rect 160343 -25462 164348 -25419
rect 160343 -25581 160369 -25462
rect 164290 -25581 164348 -25462
rect 160343 -26084 164348 -25581
rect 160343 -26118 160358 -26084
rect 164326 -26118 164348 -26084
rect 160343 -26134 164348 -26118
rect 156737 -27209 156781 -27179
rect 159452 -26494 164356 -26457
rect 159452 -26528 160358 -26494
rect 164326 -26528 164356 -26494
rect 159452 -27008 164356 -26528
rect 159452 -27054 165892 -27008
rect 159452 -27461 165785 -27054
rect 157051 -27462 165785 -27461
rect 156707 -27486 165785 -27462
rect 165855 -27486 165892 -27054
rect 156707 -27567 165892 -27486
rect 168611 -27054 168750 -27022
rect 168611 -27486 168647 -27054
rect 168717 -27486 168750 -27054
rect 156707 -27951 164356 -27567
rect 168611 -27925 168750 -27486
rect 156707 -29795 157450 -27951
rect 166918 -27962 169100 -27925
rect 166918 -28086 168798 -27962
rect 166918 -28142 166954 -28086
rect 167598 -28142 168798 -28086
rect 166918 -28180 168798 -28142
rect 169059 -28180 169100 -27962
rect 166918 -28213 169100 -28180
rect 166918 -28506 167630 -28213
rect 146808 -30684 156508 -30672
rect 146808 -30726 146820 -30684
rect 156480 -30726 156508 -30684
rect 146808 -30732 156508 -30726
rect 146802 -30748 156508 -30732
rect 157842 -30684 167562 -30674
rect 157842 -30726 157854 -30684
rect 167514 -30726 167562 -30684
rect 157842 -30748 167562 -30726
rect 146802 -30864 167562 -30748
rect 146802 -30872 157880 -30864
rect 146802 -30932 146826 -30872
rect 156448 -30924 157880 -30872
rect 167502 -30924 167562 -30864
rect 156448 -30932 167562 -30924
rect 146802 -30944 167562 -30932
rect 146802 -30952 157862 -30944
<< via1 >>
rect 156691 -27179 156752 -25046
rect 160369 -25581 164290 -25462
rect 166954 -28142 167598 -28086
rect 168798 -28180 169059 -27962
rect 146826 -30932 156448 -30872
rect 157880 -30924 167502 -30864
<< metal2 >>
rect 156671 -20621 158155 -20476
rect 156671 -21624 156772 -20621
rect 158071 -21624 158155 -20621
rect 156671 -25046 158155 -21624
rect 156671 -27179 156691 -25046
rect 156752 -27179 158155 -25046
rect 160343 -24990 164348 -24939
rect 160343 -25124 160409 -24990
rect 164292 -25124 164348 -24990
rect 160343 -25462 164348 -25124
rect 160343 -25581 160369 -25462
rect 164290 -25581 164348 -25462
rect 160343 -25604 164348 -25581
rect 156671 -27209 158155 -27179
rect 168769 -27958 169780 -27925
rect 168769 -27962 169455 -27958
rect 166901 -28086 167652 -28062
rect 166901 -28096 166954 -28086
rect 167598 -28096 167652 -28086
rect 166901 -28152 166932 -28096
rect 167618 -28152 167652 -28096
rect 166901 -28196 167652 -28152
rect 168769 -28180 168798 -27962
rect 169059 -28179 169455 -27962
rect 169749 -28179 169780 -27958
rect 169059 -28180 169780 -28179
rect 168769 -28213 169780 -28180
rect 146820 -30864 167519 -30855
rect 146820 -30872 157880 -30864
rect 146820 -30932 146826 -30872
rect 156448 -30924 157880 -30872
rect 167502 -30924 167519 -30864
rect 156448 -30932 167519 -30924
rect 146820 -31352 167519 -30932
rect 146820 -31544 146837 -31352
rect 167430 -31544 167519 -31352
rect 146820 -31558 167519 -31544
<< via2 >>
rect 156772 -21624 158071 -20621
rect 160409 -25124 164292 -24990
rect 146934 -27498 156410 -27440
rect 166932 -28142 166954 -28096
rect 166954 -28142 167598 -28096
rect 167598 -28142 167618 -28096
rect 166932 -28152 167618 -28142
rect 169455 -28179 169749 -27958
rect 146837 -31544 167430 -31352
<< metal3 >>
rect 146874 14156 156352 16000
rect 146874 1932 148562 14156
rect 154644 1932 156352 14156
rect 146874 -24694 156352 1932
rect 156671 -20596 160881 -20476
rect 156671 -20621 160165 -20596
rect 156671 -21624 156772 -20621
rect 158071 -21603 160165 -20621
rect 160775 -21603 160881 -20596
rect 158071 -21624 160881 -21603
rect 156671 -21689 160881 -21624
rect 160343 -23175 164348 -23106
rect 160343 -23326 160437 -23175
rect 164241 -23326 164348 -23175
rect 160343 -24990 164348 -23326
rect 160343 -25124 160409 -24990
rect 164292 -25124 164348 -24990
rect 160343 -25164 164348 -25124
rect 146912 -27440 156428 -27432
rect 146912 -27498 146934 -27440
rect 156410 -27498 156428 -27440
rect 146912 -28138 156428 -27498
rect 169409 -27958 170803 -27925
rect 166710 -28096 167694 -28012
rect 166710 -28152 166932 -28096
rect 167618 -28152 167694 -28096
rect 166710 -28165 167694 -28152
rect 166772 -28168 167694 -28165
rect 166804 -28208 167656 -28168
rect 169409 -28179 169455 -27958
rect 169749 -27961 170803 -27958
rect 169749 -28179 170460 -27961
rect 169409 -28186 170460 -28179
rect 170764 -28186 170803 -27961
rect 169409 -28213 170803 -28186
rect 146772 -31312 168651 -31277
rect 146772 -31352 168147 -31312
rect 146772 -31544 146837 -31352
rect 167430 -31544 168147 -31352
rect 146772 -31579 168147 -31544
rect 168605 -31579 168651 -31312
rect 146772 -31615 168651 -31579
<< via3 >>
rect 148562 1932 154644 14156
rect 160165 -21603 160775 -20596
rect 160437 -23326 164241 -23175
rect 170460 -28186 170764 -27961
rect 168147 -31579 168605 -31312
<< metal4 >>
rect 159000 374980 351997 379374
rect 159000 350084 317582 374980
rect 339915 350084 351997 374980
rect 159000 344551 351997 350084
rect 146874 14932 156352 16000
rect 146874 1038 147788 14932
rect 155360 1038 156352 14932
rect 146874 0 156352 1038
rect 160074 -20549 164284 -20476
rect 160074 -20596 163186 -20549
rect 160074 -21603 160165 -20596
rect 160775 -21603 163186 -20596
rect 160074 -21645 163186 -21603
rect 163747 -21645 164284 -20549
rect 160074 -21689 164284 -21645
rect 160343 -22553 165003 -22504
rect 160343 -23175 164630 -22553
rect 160343 -23326 160437 -23175
rect 164241 -23326 164630 -23175
rect 160343 -23332 164630 -23326
rect 164903 -23332 165003 -22553
rect 160343 -23370 165003 -23332
rect 170438 -27961 171909 -27925
rect 170438 -28186 170460 -27961
rect 170764 -28186 171523 -27961
rect 170438 -28203 171523 -28186
rect 171878 -28203 171909 -27961
rect 170438 -28213 171909 -28203
rect 168109 -30786 170325 -30630
rect 168109 -31312 169819 -30786
rect 168109 -31579 168147 -31312
rect 168605 -31535 169819 -31312
rect 170140 -31535 170325 -30786
rect 168605 -31579 170325 -31535
rect 168109 -31651 170325 -31579
<< via4 >>
rect 317582 350084 339915 374980
rect 147788 14156 155360 14932
rect 147788 1932 148562 14156
rect 148562 1932 154644 14156
rect 154644 1932 155360 14156
rect 147788 1038 155360 1932
rect 163186 -21645 163747 -20549
rect 164630 -23332 164903 -22553
rect 171523 -28203 171878 -27961
rect 169819 -31535 170140 -30786
<< metal5 >>
rect 313801 374980 352952 379374
rect 313801 350084 317582 374980
rect 339915 350084 352952 374980
rect 313801 344551 352952 350084
rect 146874 14932 156352 16000
rect 146874 1038 147788 14932
rect 155360 1038 156352 14932
rect 146874 0 156352 1038
rect 163107 -20549 167317 -20476
rect 163107 -21645 163186 -20549
rect 163747 -21645 167317 -20549
rect 163107 -21689 167317 -21645
rect 164597 -22553 169257 -22504
rect 164597 -23332 164630 -22553
rect 164903 -23332 169257 -22553
rect 164597 -23370 169257 -23332
rect 171445 -27961 172056 -27810
rect 171445 -28203 171523 -27961
rect 171878 -28203 172056 -27961
rect 171445 -28303 172056 -28203
rect 169750 -30786 171581 -30396
rect 169750 -31535 169819 -30786
rect 170140 -31535 171581 -30786
rect 169750 -31847 171581 -31535
use sky130_fd_pr__res_generic_po_u1tz6h  sky130_fd_pr__res_generic_po_u1tz6h_0
timestamp 1606531739
transform 1 0 162342 0 1 -26306
box -2166 -404 2166 404
use sky130_fd_pr__res_high_po_0p35_i8je6j  sky130_fd_pr__res_high_po_0p35_i8je6j_0
timestamp 1606531739
transform 1 0 167251 0 1 -26054
box -1632 -1598 1632 1598
use transistor_1m  transistor_1m_2
timestamp 1606422944
transform 1 0 128835 0 1 -31687
box 28887 745 38986 3606
use transistor_1m  transistor_1m_1
timestamp 1606422944
transform 1 0 117795 0 1 -31685
box 28887 745 38986 3606
use transistor_1m  transistor_1m_0
timestamp 1606422944
transform 1 0 117759 0 1 -28251
box 28887 745 38986 3606
use INDUCTOR_L  INDUCTOR_L_0
timestamp 1606452767
transform 1 0 432600 0 1 171000
box -432600 -171000 -79800 178200
<< labels >>
rlabel metal5 342989 346603 346877 377149 1 vdd
port 1 n
rlabel metal5 166668 -21526 167008 -20656 1 Vgate
port 2 n
rlabel metal5 171926 -28261 172027 -27853 1 Isource
port 3 n
rlabel metal5 168834 -23282 169169 -22611 1 Rnode
port 4 n
rlabel metal5 171123 -31584 171405 -30698 1 vss
port 5 n
rlabel metal3 147547 -13778 155259 -3811 1 out
<< end >>
