magic
tech sky130A
magscale 1 2
timestamp 1606471058
<< pwell >>
rect -2457 -910 2457 910
<< nmoslvt >>
rect -2261 -700 -1861 700
rect -1803 -700 -1403 700
rect -1345 -700 -945 700
rect -887 -700 -487 700
rect -429 -700 -29 700
rect 29 -700 429 700
rect 487 -700 887 700
rect 945 -700 1345 700
rect 1403 -700 1803 700
rect 1861 -700 2261 700
<< ndiff >>
rect -2319 688 -2261 700
rect -2319 -688 -2307 688
rect -2273 -688 -2261 688
rect -2319 -700 -2261 -688
rect -1861 688 -1803 700
rect -1861 -688 -1849 688
rect -1815 -688 -1803 688
rect -1861 -700 -1803 -688
rect -1403 688 -1345 700
rect -1403 -688 -1391 688
rect -1357 -688 -1345 688
rect -1403 -700 -1345 -688
rect -945 688 -887 700
rect -945 -688 -933 688
rect -899 -688 -887 688
rect -945 -700 -887 -688
rect -487 688 -429 700
rect -487 -688 -475 688
rect -441 -688 -429 688
rect -487 -700 -429 -688
rect -29 688 29 700
rect -29 -688 -17 688
rect 17 -688 29 688
rect -29 -700 29 -688
rect 429 688 487 700
rect 429 -688 441 688
rect 475 -688 487 688
rect 429 -700 487 -688
rect 887 688 945 700
rect 887 -688 899 688
rect 933 -688 945 688
rect 887 -700 945 -688
rect 1345 688 1403 700
rect 1345 -688 1357 688
rect 1391 -688 1403 688
rect 1345 -700 1403 -688
rect 1803 688 1861 700
rect 1803 -688 1815 688
rect 1849 -688 1861 688
rect 1803 -700 1861 -688
rect 2261 688 2319 700
rect 2261 -688 2273 688
rect 2307 -688 2319 688
rect 2261 -700 2319 -688
<< ndiffc >>
rect -2307 -688 -2273 688
rect -1849 -688 -1815 688
rect -1391 -688 -1357 688
rect -933 -688 -899 688
rect -475 -688 -441 688
rect -17 -688 17 688
rect 441 -688 475 688
rect 899 -688 933 688
rect 1357 -688 1391 688
rect 1815 -688 1849 688
rect 2273 -688 2307 688
<< psubdiff >>
rect -2421 840 -2325 874
rect 2325 840 2421 874
rect -2421 778 -2387 840
rect 2387 778 2421 840
rect -2421 -840 -2387 -778
rect 2387 -840 2421 -778
rect -2421 -874 -2325 -840
rect 2325 -874 2421 -840
<< psubdiffcont >>
rect -2325 840 2325 874
rect -2421 -778 -2387 778
rect 2387 -778 2421 778
rect -2325 -874 2325 -840
<< poly >>
rect -2261 772 -1861 788
rect -2261 738 -2245 772
rect -1877 738 -1861 772
rect -2261 700 -1861 738
rect -1803 772 -1403 788
rect -1803 738 -1787 772
rect -1419 738 -1403 772
rect -1803 700 -1403 738
rect -1345 772 -945 788
rect -1345 738 -1329 772
rect -961 738 -945 772
rect -1345 700 -945 738
rect -887 772 -487 788
rect -887 738 -871 772
rect -503 738 -487 772
rect -887 700 -487 738
rect -429 772 -29 788
rect -429 738 -413 772
rect -45 738 -29 772
rect -429 700 -29 738
rect 29 772 429 788
rect 29 738 45 772
rect 413 738 429 772
rect 29 700 429 738
rect 487 772 887 788
rect 487 738 503 772
rect 871 738 887 772
rect 487 700 887 738
rect 945 772 1345 788
rect 945 738 961 772
rect 1329 738 1345 772
rect 945 700 1345 738
rect 1403 772 1803 788
rect 1403 738 1419 772
rect 1787 738 1803 772
rect 1403 700 1803 738
rect 1861 772 2261 788
rect 1861 738 1877 772
rect 2245 738 2261 772
rect 1861 700 2261 738
rect -2261 -738 -1861 -700
rect -2261 -772 -2245 -738
rect -1877 -772 -1861 -738
rect -2261 -788 -1861 -772
rect -1803 -738 -1403 -700
rect -1803 -772 -1787 -738
rect -1419 -772 -1403 -738
rect -1803 -788 -1403 -772
rect -1345 -738 -945 -700
rect -1345 -772 -1329 -738
rect -961 -772 -945 -738
rect -1345 -788 -945 -772
rect -887 -738 -487 -700
rect -887 -772 -871 -738
rect -503 -772 -487 -738
rect -887 -788 -487 -772
rect -429 -738 -29 -700
rect -429 -772 -413 -738
rect -45 -772 -29 -738
rect -429 -788 -29 -772
rect 29 -738 429 -700
rect 29 -772 45 -738
rect 413 -772 429 -738
rect 29 -788 429 -772
rect 487 -738 887 -700
rect 487 -772 503 -738
rect 871 -772 887 -738
rect 487 -788 887 -772
rect 945 -738 1345 -700
rect 945 -772 961 -738
rect 1329 -772 1345 -738
rect 945 -788 1345 -772
rect 1403 -738 1803 -700
rect 1403 -772 1419 -738
rect 1787 -772 1803 -738
rect 1403 -788 1803 -772
rect 1861 -738 2261 -700
rect 1861 -772 1877 -738
rect 2245 -772 2261 -738
rect 1861 -788 2261 -772
<< polycont >>
rect -2245 738 -1877 772
rect -1787 738 -1419 772
rect -1329 738 -961 772
rect -871 738 -503 772
rect -413 738 -45 772
rect 45 738 413 772
rect 503 738 871 772
rect 961 738 1329 772
rect 1419 738 1787 772
rect 1877 738 2245 772
rect -2245 -772 -1877 -738
rect -1787 -772 -1419 -738
rect -1329 -772 -961 -738
rect -871 -772 -503 -738
rect -413 -772 -45 -738
rect 45 -772 413 -738
rect 503 -772 871 -738
rect 961 -772 1329 -738
rect 1419 -772 1787 -738
rect 1877 -772 2245 -738
<< locali >>
rect -2421 840 -2325 874
rect 2325 840 2421 874
rect -2421 778 -2387 840
rect 2387 778 2421 840
rect -2261 738 -2245 772
rect -1877 738 -1861 772
rect -1803 738 -1787 772
rect -1419 738 -1403 772
rect -1345 738 -1329 772
rect -961 738 -945 772
rect -887 738 -871 772
rect -503 738 -487 772
rect -429 738 -413 772
rect -45 738 -29 772
rect 29 738 45 772
rect 413 738 429 772
rect 487 738 503 772
rect 871 738 887 772
rect 945 738 961 772
rect 1329 738 1345 772
rect 1403 738 1419 772
rect 1787 738 1803 772
rect 1861 738 1877 772
rect 2245 738 2261 772
rect -2307 688 -2273 704
rect -2307 -704 -2273 -688
rect -1849 688 -1815 704
rect -1849 -704 -1815 -688
rect -1391 688 -1357 704
rect -1391 -704 -1357 -688
rect -933 688 -899 704
rect -933 -704 -899 -688
rect -475 688 -441 704
rect -475 -704 -441 -688
rect -17 688 17 704
rect -17 -704 17 -688
rect 441 688 475 704
rect 441 -704 475 -688
rect 899 688 933 704
rect 899 -704 933 -688
rect 1357 688 1391 704
rect 1357 -704 1391 -688
rect 1815 688 1849 704
rect 1815 -704 1849 -688
rect 2273 688 2307 704
rect 2273 -704 2307 -688
rect -2261 -772 -2245 -738
rect -1877 -772 -1861 -738
rect -1803 -772 -1787 -738
rect -1419 -772 -1403 -738
rect -1345 -772 -1329 -738
rect -961 -772 -945 -738
rect -887 -772 -871 -738
rect -503 -772 -487 -738
rect -429 -772 -413 -738
rect -45 -772 -29 -738
rect 29 -772 45 -738
rect 413 -772 429 -738
rect 487 -772 503 -738
rect 871 -772 887 -738
rect 945 -772 961 -738
rect 1329 -772 1345 -738
rect 1403 -772 1419 -738
rect 1787 -772 1803 -738
rect 1861 -772 1877 -738
rect 2245 -772 2261 -738
rect -2421 -840 -2387 -778
rect 2387 -840 2421 -778
rect -2421 -874 -2325 -840
rect 2325 -874 2421 -840
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -2404 -857 2404 857
string parameters w 7 l 2 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
