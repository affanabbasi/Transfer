magic
tech sky130A
magscale 1 2
timestamp 1606421359
<< pwell >>
rect -4967 -1210 4967 1210
<< nmos >>
rect -4767 -1000 -4737 1000
rect -4671 -1000 -4641 1000
rect -4575 -1000 -4545 1000
rect -4479 -1000 -4449 1000
rect -4383 -1000 -4353 1000
rect -4287 -1000 -4257 1000
rect -4191 -1000 -4161 1000
rect -4095 -1000 -4065 1000
rect -3999 -1000 -3969 1000
rect -3903 -1000 -3873 1000
rect -3807 -1000 -3777 1000
rect -3711 -1000 -3681 1000
rect -3615 -1000 -3585 1000
rect -3519 -1000 -3489 1000
rect -3423 -1000 -3393 1000
rect -3327 -1000 -3297 1000
rect -3231 -1000 -3201 1000
rect -3135 -1000 -3105 1000
rect -3039 -1000 -3009 1000
rect -2943 -1000 -2913 1000
rect -2847 -1000 -2817 1000
rect -2751 -1000 -2721 1000
rect -2655 -1000 -2625 1000
rect -2559 -1000 -2529 1000
rect -2463 -1000 -2433 1000
rect -2367 -1000 -2337 1000
rect -2271 -1000 -2241 1000
rect -2175 -1000 -2145 1000
rect -2079 -1000 -2049 1000
rect -1983 -1000 -1953 1000
rect -1887 -1000 -1857 1000
rect -1791 -1000 -1761 1000
rect -1695 -1000 -1665 1000
rect -1599 -1000 -1569 1000
rect -1503 -1000 -1473 1000
rect -1407 -1000 -1377 1000
rect -1311 -1000 -1281 1000
rect -1215 -1000 -1185 1000
rect -1119 -1000 -1089 1000
rect -1023 -1000 -993 1000
rect -927 -1000 -897 1000
rect -831 -1000 -801 1000
rect -735 -1000 -705 1000
rect -639 -1000 -609 1000
rect -543 -1000 -513 1000
rect -447 -1000 -417 1000
rect -351 -1000 -321 1000
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
rect 321 -1000 351 1000
rect 417 -1000 447 1000
rect 513 -1000 543 1000
rect 609 -1000 639 1000
rect 705 -1000 735 1000
rect 801 -1000 831 1000
rect 897 -1000 927 1000
rect 993 -1000 1023 1000
rect 1089 -1000 1119 1000
rect 1185 -1000 1215 1000
rect 1281 -1000 1311 1000
rect 1377 -1000 1407 1000
rect 1473 -1000 1503 1000
rect 1569 -1000 1599 1000
rect 1665 -1000 1695 1000
rect 1761 -1000 1791 1000
rect 1857 -1000 1887 1000
rect 1953 -1000 1983 1000
rect 2049 -1000 2079 1000
rect 2145 -1000 2175 1000
rect 2241 -1000 2271 1000
rect 2337 -1000 2367 1000
rect 2433 -1000 2463 1000
rect 2529 -1000 2559 1000
rect 2625 -1000 2655 1000
rect 2721 -1000 2751 1000
rect 2817 -1000 2847 1000
rect 2913 -1000 2943 1000
rect 3009 -1000 3039 1000
rect 3105 -1000 3135 1000
rect 3201 -1000 3231 1000
rect 3297 -1000 3327 1000
rect 3393 -1000 3423 1000
rect 3489 -1000 3519 1000
rect 3585 -1000 3615 1000
rect 3681 -1000 3711 1000
rect 3777 -1000 3807 1000
rect 3873 -1000 3903 1000
rect 3969 -1000 3999 1000
rect 4065 -1000 4095 1000
rect 4161 -1000 4191 1000
rect 4257 -1000 4287 1000
rect 4353 -1000 4383 1000
rect 4449 -1000 4479 1000
rect 4545 -1000 4575 1000
rect 4641 -1000 4671 1000
rect 4737 -1000 4767 1000
<< ndiff >>
rect -4829 988 -4767 1000
rect -4829 -988 -4817 988
rect -4783 -988 -4767 988
rect -4829 -1000 -4767 -988
rect -4737 988 -4671 1000
rect -4737 -988 -4721 988
rect -4687 -988 -4671 988
rect -4737 -1000 -4671 -988
rect -4641 988 -4575 1000
rect -4641 -988 -4625 988
rect -4591 -988 -4575 988
rect -4641 -1000 -4575 -988
rect -4545 988 -4479 1000
rect -4545 -988 -4529 988
rect -4495 -988 -4479 988
rect -4545 -1000 -4479 -988
rect -4449 988 -4383 1000
rect -4449 -988 -4433 988
rect -4399 -988 -4383 988
rect -4449 -1000 -4383 -988
rect -4353 988 -4287 1000
rect -4353 -988 -4337 988
rect -4303 -988 -4287 988
rect -4353 -1000 -4287 -988
rect -4257 988 -4191 1000
rect -4257 -988 -4241 988
rect -4207 -988 -4191 988
rect -4257 -1000 -4191 -988
rect -4161 988 -4095 1000
rect -4161 -988 -4145 988
rect -4111 -988 -4095 988
rect -4161 -1000 -4095 -988
rect -4065 988 -3999 1000
rect -4065 -988 -4049 988
rect -4015 -988 -3999 988
rect -4065 -1000 -3999 -988
rect -3969 988 -3903 1000
rect -3969 -988 -3953 988
rect -3919 -988 -3903 988
rect -3969 -1000 -3903 -988
rect -3873 988 -3807 1000
rect -3873 -988 -3857 988
rect -3823 -988 -3807 988
rect -3873 -1000 -3807 -988
rect -3777 988 -3711 1000
rect -3777 -988 -3761 988
rect -3727 -988 -3711 988
rect -3777 -1000 -3711 -988
rect -3681 988 -3615 1000
rect -3681 -988 -3665 988
rect -3631 -988 -3615 988
rect -3681 -1000 -3615 -988
rect -3585 988 -3519 1000
rect -3585 -988 -3569 988
rect -3535 -988 -3519 988
rect -3585 -1000 -3519 -988
rect -3489 988 -3423 1000
rect -3489 -988 -3473 988
rect -3439 -988 -3423 988
rect -3489 -1000 -3423 -988
rect -3393 988 -3327 1000
rect -3393 -988 -3377 988
rect -3343 -988 -3327 988
rect -3393 -1000 -3327 -988
rect -3297 988 -3231 1000
rect -3297 -988 -3281 988
rect -3247 -988 -3231 988
rect -3297 -1000 -3231 -988
rect -3201 988 -3135 1000
rect -3201 -988 -3185 988
rect -3151 -988 -3135 988
rect -3201 -1000 -3135 -988
rect -3105 988 -3039 1000
rect -3105 -988 -3089 988
rect -3055 -988 -3039 988
rect -3105 -1000 -3039 -988
rect -3009 988 -2943 1000
rect -3009 -988 -2993 988
rect -2959 -988 -2943 988
rect -3009 -1000 -2943 -988
rect -2913 988 -2847 1000
rect -2913 -988 -2897 988
rect -2863 -988 -2847 988
rect -2913 -1000 -2847 -988
rect -2817 988 -2751 1000
rect -2817 -988 -2801 988
rect -2767 -988 -2751 988
rect -2817 -1000 -2751 -988
rect -2721 988 -2655 1000
rect -2721 -988 -2705 988
rect -2671 -988 -2655 988
rect -2721 -1000 -2655 -988
rect -2625 988 -2559 1000
rect -2625 -988 -2609 988
rect -2575 -988 -2559 988
rect -2625 -1000 -2559 -988
rect -2529 988 -2463 1000
rect -2529 -988 -2513 988
rect -2479 -988 -2463 988
rect -2529 -1000 -2463 -988
rect -2433 988 -2367 1000
rect -2433 -988 -2417 988
rect -2383 -988 -2367 988
rect -2433 -1000 -2367 -988
rect -2337 988 -2271 1000
rect -2337 -988 -2321 988
rect -2287 -988 -2271 988
rect -2337 -1000 -2271 -988
rect -2241 988 -2175 1000
rect -2241 -988 -2225 988
rect -2191 -988 -2175 988
rect -2241 -1000 -2175 -988
rect -2145 988 -2079 1000
rect -2145 -988 -2129 988
rect -2095 -988 -2079 988
rect -2145 -1000 -2079 -988
rect -2049 988 -1983 1000
rect -2049 -988 -2033 988
rect -1999 -988 -1983 988
rect -2049 -1000 -1983 -988
rect -1953 988 -1887 1000
rect -1953 -988 -1937 988
rect -1903 -988 -1887 988
rect -1953 -1000 -1887 -988
rect -1857 988 -1791 1000
rect -1857 -988 -1841 988
rect -1807 -988 -1791 988
rect -1857 -1000 -1791 -988
rect -1761 988 -1695 1000
rect -1761 -988 -1745 988
rect -1711 -988 -1695 988
rect -1761 -1000 -1695 -988
rect -1665 988 -1599 1000
rect -1665 -988 -1649 988
rect -1615 -988 -1599 988
rect -1665 -1000 -1599 -988
rect -1569 988 -1503 1000
rect -1569 -988 -1553 988
rect -1519 -988 -1503 988
rect -1569 -1000 -1503 -988
rect -1473 988 -1407 1000
rect -1473 -988 -1457 988
rect -1423 -988 -1407 988
rect -1473 -1000 -1407 -988
rect -1377 988 -1311 1000
rect -1377 -988 -1361 988
rect -1327 -988 -1311 988
rect -1377 -1000 -1311 -988
rect -1281 988 -1215 1000
rect -1281 -988 -1265 988
rect -1231 -988 -1215 988
rect -1281 -1000 -1215 -988
rect -1185 988 -1119 1000
rect -1185 -988 -1169 988
rect -1135 -988 -1119 988
rect -1185 -1000 -1119 -988
rect -1089 988 -1023 1000
rect -1089 -988 -1073 988
rect -1039 -988 -1023 988
rect -1089 -1000 -1023 -988
rect -993 988 -927 1000
rect -993 -988 -977 988
rect -943 -988 -927 988
rect -993 -1000 -927 -988
rect -897 988 -831 1000
rect -897 -988 -881 988
rect -847 -988 -831 988
rect -897 -1000 -831 -988
rect -801 988 -735 1000
rect -801 -988 -785 988
rect -751 -988 -735 988
rect -801 -1000 -735 -988
rect -705 988 -639 1000
rect -705 -988 -689 988
rect -655 -988 -639 988
rect -705 -1000 -639 -988
rect -609 988 -543 1000
rect -609 -988 -593 988
rect -559 -988 -543 988
rect -609 -1000 -543 -988
rect -513 988 -447 1000
rect -513 -988 -497 988
rect -463 -988 -447 988
rect -513 -1000 -447 -988
rect -417 988 -351 1000
rect -417 -988 -401 988
rect -367 -988 -351 988
rect -417 -1000 -351 -988
rect -321 988 -255 1000
rect -321 -988 -305 988
rect -271 -988 -255 988
rect -321 -1000 -255 -988
rect -225 988 -159 1000
rect -225 -988 -209 988
rect -175 -988 -159 988
rect -225 -1000 -159 -988
rect -129 988 -63 1000
rect -129 -988 -113 988
rect -79 -988 -63 988
rect -129 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 129 1000
rect 63 -988 79 988
rect 113 -988 129 988
rect 63 -1000 129 -988
rect 159 988 225 1000
rect 159 -988 175 988
rect 209 -988 225 988
rect 159 -1000 225 -988
rect 255 988 321 1000
rect 255 -988 271 988
rect 305 -988 321 988
rect 255 -1000 321 -988
rect 351 988 417 1000
rect 351 -988 367 988
rect 401 -988 417 988
rect 351 -1000 417 -988
rect 447 988 513 1000
rect 447 -988 463 988
rect 497 -988 513 988
rect 447 -1000 513 -988
rect 543 988 609 1000
rect 543 -988 559 988
rect 593 -988 609 988
rect 543 -1000 609 -988
rect 639 988 705 1000
rect 639 -988 655 988
rect 689 -988 705 988
rect 639 -1000 705 -988
rect 735 988 801 1000
rect 735 -988 751 988
rect 785 -988 801 988
rect 735 -1000 801 -988
rect 831 988 897 1000
rect 831 -988 847 988
rect 881 -988 897 988
rect 831 -1000 897 -988
rect 927 988 993 1000
rect 927 -988 943 988
rect 977 -988 993 988
rect 927 -1000 993 -988
rect 1023 988 1089 1000
rect 1023 -988 1039 988
rect 1073 -988 1089 988
rect 1023 -1000 1089 -988
rect 1119 988 1185 1000
rect 1119 -988 1135 988
rect 1169 -988 1185 988
rect 1119 -1000 1185 -988
rect 1215 988 1281 1000
rect 1215 -988 1231 988
rect 1265 -988 1281 988
rect 1215 -1000 1281 -988
rect 1311 988 1377 1000
rect 1311 -988 1327 988
rect 1361 -988 1377 988
rect 1311 -1000 1377 -988
rect 1407 988 1473 1000
rect 1407 -988 1423 988
rect 1457 -988 1473 988
rect 1407 -1000 1473 -988
rect 1503 988 1569 1000
rect 1503 -988 1519 988
rect 1553 -988 1569 988
rect 1503 -1000 1569 -988
rect 1599 988 1665 1000
rect 1599 -988 1615 988
rect 1649 -988 1665 988
rect 1599 -1000 1665 -988
rect 1695 988 1761 1000
rect 1695 -988 1711 988
rect 1745 -988 1761 988
rect 1695 -1000 1761 -988
rect 1791 988 1857 1000
rect 1791 -988 1807 988
rect 1841 -988 1857 988
rect 1791 -1000 1857 -988
rect 1887 988 1953 1000
rect 1887 -988 1903 988
rect 1937 -988 1953 988
rect 1887 -1000 1953 -988
rect 1983 988 2049 1000
rect 1983 -988 1999 988
rect 2033 -988 2049 988
rect 1983 -1000 2049 -988
rect 2079 988 2145 1000
rect 2079 -988 2095 988
rect 2129 -988 2145 988
rect 2079 -1000 2145 -988
rect 2175 988 2241 1000
rect 2175 -988 2191 988
rect 2225 -988 2241 988
rect 2175 -1000 2241 -988
rect 2271 988 2337 1000
rect 2271 -988 2287 988
rect 2321 -988 2337 988
rect 2271 -1000 2337 -988
rect 2367 988 2433 1000
rect 2367 -988 2383 988
rect 2417 -988 2433 988
rect 2367 -1000 2433 -988
rect 2463 988 2529 1000
rect 2463 -988 2479 988
rect 2513 -988 2529 988
rect 2463 -1000 2529 -988
rect 2559 988 2625 1000
rect 2559 -988 2575 988
rect 2609 -988 2625 988
rect 2559 -1000 2625 -988
rect 2655 988 2721 1000
rect 2655 -988 2671 988
rect 2705 -988 2721 988
rect 2655 -1000 2721 -988
rect 2751 988 2817 1000
rect 2751 -988 2767 988
rect 2801 -988 2817 988
rect 2751 -1000 2817 -988
rect 2847 988 2913 1000
rect 2847 -988 2863 988
rect 2897 -988 2913 988
rect 2847 -1000 2913 -988
rect 2943 988 3009 1000
rect 2943 -988 2959 988
rect 2993 -988 3009 988
rect 2943 -1000 3009 -988
rect 3039 988 3105 1000
rect 3039 -988 3055 988
rect 3089 -988 3105 988
rect 3039 -1000 3105 -988
rect 3135 988 3201 1000
rect 3135 -988 3151 988
rect 3185 -988 3201 988
rect 3135 -1000 3201 -988
rect 3231 988 3297 1000
rect 3231 -988 3247 988
rect 3281 -988 3297 988
rect 3231 -1000 3297 -988
rect 3327 988 3393 1000
rect 3327 -988 3343 988
rect 3377 -988 3393 988
rect 3327 -1000 3393 -988
rect 3423 988 3489 1000
rect 3423 -988 3439 988
rect 3473 -988 3489 988
rect 3423 -1000 3489 -988
rect 3519 988 3585 1000
rect 3519 -988 3535 988
rect 3569 -988 3585 988
rect 3519 -1000 3585 -988
rect 3615 988 3681 1000
rect 3615 -988 3631 988
rect 3665 -988 3681 988
rect 3615 -1000 3681 -988
rect 3711 988 3777 1000
rect 3711 -988 3727 988
rect 3761 -988 3777 988
rect 3711 -1000 3777 -988
rect 3807 988 3873 1000
rect 3807 -988 3823 988
rect 3857 -988 3873 988
rect 3807 -1000 3873 -988
rect 3903 988 3969 1000
rect 3903 -988 3919 988
rect 3953 -988 3969 988
rect 3903 -1000 3969 -988
rect 3999 988 4065 1000
rect 3999 -988 4015 988
rect 4049 -988 4065 988
rect 3999 -1000 4065 -988
rect 4095 988 4161 1000
rect 4095 -988 4111 988
rect 4145 -988 4161 988
rect 4095 -1000 4161 -988
rect 4191 988 4257 1000
rect 4191 -988 4207 988
rect 4241 -988 4257 988
rect 4191 -1000 4257 -988
rect 4287 988 4353 1000
rect 4287 -988 4303 988
rect 4337 -988 4353 988
rect 4287 -1000 4353 -988
rect 4383 988 4449 1000
rect 4383 -988 4399 988
rect 4433 -988 4449 988
rect 4383 -1000 4449 -988
rect 4479 988 4545 1000
rect 4479 -988 4495 988
rect 4529 -988 4545 988
rect 4479 -1000 4545 -988
rect 4575 988 4641 1000
rect 4575 -988 4591 988
rect 4625 -988 4641 988
rect 4575 -1000 4641 -988
rect 4671 988 4737 1000
rect 4671 -988 4687 988
rect 4721 -988 4737 988
rect 4671 -1000 4737 -988
rect 4767 988 4829 1000
rect 4767 -988 4783 988
rect 4817 -988 4829 988
rect 4767 -1000 4829 -988
<< ndiffc >>
rect -4817 -988 -4783 988
rect -4721 -988 -4687 988
rect -4625 -988 -4591 988
rect -4529 -988 -4495 988
rect -4433 -988 -4399 988
rect -4337 -988 -4303 988
rect -4241 -988 -4207 988
rect -4145 -988 -4111 988
rect -4049 -988 -4015 988
rect -3953 -988 -3919 988
rect -3857 -988 -3823 988
rect -3761 -988 -3727 988
rect -3665 -988 -3631 988
rect -3569 -988 -3535 988
rect -3473 -988 -3439 988
rect -3377 -988 -3343 988
rect -3281 -988 -3247 988
rect -3185 -988 -3151 988
rect -3089 -988 -3055 988
rect -2993 -988 -2959 988
rect -2897 -988 -2863 988
rect -2801 -988 -2767 988
rect -2705 -988 -2671 988
rect -2609 -988 -2575 988
rect -2513 -988 -2479 988
rect -2417 -988 -2383 988
rect -2321 -988 -2287 988
rect -2225 -988 -2191 988
rect -2129 -988 -2095 988
rect -2033 -988 -1999 988
rect -1937 -988 -1903 988
rect -1841 -988 -1807 988
rect -1745 -988 -1711 988
rect -1649 -988 -1615 988
rect -1553 -988 -1519 988
rect -1457 -988 -1423 988
rect -1361 -988 -1327 988
rect -1265 -988 -1231 988
rect -1169 -988 -1135 988
rect -1073 -988 -1039 988
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect 1039 -988 1073 988
rect 1135 -988 1169 988
rect 1231 -988 1265 988
rect 1327 -988 1361 988
rect 1423 -988 1457 988
rect 1519 -988 1553 988
rect 1615 -988 1649 988
rect 1711 -988 1745 988
rect 1807 -988 1841 988
rect 1903 -988 1937 988
rect 1999 -988 2033 988
rect 2095 -988 2129 988
rect 2191 -988 2225 988
rect 2287 -988 2321 988
rect 2383 -988 2417 988
rect 2479 -988 2513 988
rect 2575 -988 2609 988
rect 2671 -988 2705 988
rect 2767 -988 2801 988
rect 2863 -988 2897 988
rect 2959 -988 2993 988
rect 3055 -988 3089 988
rect 3151 -988 3185 988
rect 3247 -988 3281 988
rect 3343 -988 3377 988
rect 3439 -988 3473 988
rect 3535 -988 3569 988
rect 3631 -988 3665 988
rect 3727 -988 3761 988
rect 3823 -988 3857 988
rect 3919 -988 3953 988
rect 4015 -988 4049 988
rect 4111 -988 4145 988
rect 4207 -988 4241 988
rect 4303 -988 4337 988
rect 4399 -988 4433 988
rect 4495 -988 4529 988
rect 4591 -988 4625 988
rect 4687 -988 4721 988
rect 4783 -988 4817 988
<< psubdiff >>
rect -4931 1140 -4835 1174
rect 4835 1140 4931 1174
rect -4931 1078 -4897 1140
rect 4897 1078 4931 1140
rect -4931 -1140 -4897 -1078
rect 4897 -1140 4931 -1078
rect -4931 -1174 -4835 -1140
rect 4835 -1174 4931 -1140
<< psubdiffcont >>
rect -4835 1140 4835 1174
rect -4931 -1078 -4897 1078
rect 4897 -1078 4931 1078
rect -4835 -1174 4835 -1140
<< poly >>
rect -4689 1072 -4623 1088
rect -4689 1038 -4673 1072
rect -4639 1038 -4623 1072
rect -4767 1000 -4737 1026
rect -4689 1022 -4623 1038
rect -4497 1072 -4431 1088
rect -4497 1038 -4481 1072
rect -4447 1038 -4431 1072
rect -4671 1000 -4641 1022
rect -4575 1000 -4545 1026
rect -4497 1022 -4431 1038
rect -4305 1072 -4239 1088
rect -4305 1038 -4289 1072
rect -4255 1038 -4239 1072
rect -4479 1000 -4449 1022
rect -4383 1000 -4353 1026
rect -4305 1022 -4239 1038
rect -4113 1072 -4047 1088
rect -4113 1038 -4097 1072
rect -4063 1038 -4047 1072
rect -4287 1000 -4257 1022
rect -4191 1000 -4161 1026
rect -4113 1022 -4047 1038
rect -3921 1072 -3855 1088
rect -3921 1038 -3905 1072
rect -3871 1038 -3855 1072
rect -4095 1000 -4065 1022
rect -3999 1000 -3969 1026
rect -3921 1022 -3855 1038
rect -3729 1072 -3663 1088
rect -3729 1038 -3713 1072
rect -3679 1038 -3663 1072
rect -3903 1000 -3873 1022
rect -3807 1000 -3777 1026
rect -3729 1022 -3663 1038
rect -3537 1072 -3471 1088
rect -3537 1038 -3521 1072
rect -3487 1038 -3471 1072
rect -3711 1000 -3681 1022
rect -3615 1000 -3585 1026
rect -3537 1022 -3471 1038
rect -3345 1072 -3279 1088
rect -3345 1038 -3329 1072
rect -3295 1038 -3279 1072
rect -3519 1000 -3489 1022
rect -3423 1000 -3393 1026
rect -3345 1022 -3279 1038
rect -3153 1072 -3087 1088
rect -3153 1038 -3137 1072
rect -3103 1038 -3087 1072
rect -3327 1000 -3297 1022
rect -3231 1000 -3201 1026
rect -3153 1022 -3087 1038
rect -2961 1072 -2895 1088
rect -2961 1038 -2945 1072
rect -2911 1038 -2895 1072
rect -3135 1000 -3105 1022
rect -3039 1000 -3009 1026
rect -2961 1022 -2895 1038
rect -2769 1072 -2703 1088
rect -2769 1038 -2753 1072
rect -2719 1038 -2703 1072
rect -2943 1000 -2913 1022
rect -2847 1000 -2817 1026
rect -2769 1022 -2703 1038
rect -2577 1072 -2511 1088
rect -2577 1038 -2561 1072
rect -2527 1038 -2511 1072
rect -2751 1000 -2721 1022
rect -2655 1000 -2625 1026
rect -2577 1022 -2511 1038
rect -2385 1072 -2319 1088
rect -2385 1038 -2369 1072
rect -2335 1038 -2319 1072
rect -2559 1000 -2529 1022
rect -2463 1000 -2433 1026
rect -2385 1022 -2319 1038
rect -2193 1072 -2127 1088
rect -2193 1038 -2177 1072
rect -2143 1038 -2127 1072
rect -2367 1000 -2337 1022
rect -2271 1000 -2241 1026
rect -2193 1022 -2127 1038
rect -2001 1072 -1935 1088
rect -2001 1038 -1985 1072
rect -1951 1038 -1935 1072
rect -2175 1000 -2145 1022
rect -2079 1000 -2049 1026
rect -2001 1022 -1935 1038
rect -1809 1072 -1743 1088
rect -1809 1038 -1793 1072
rect -1759 1038 -1743 1072
rect -1983 1000 -1953 1022
rect -1887 1000 -1857 1026
rect -1809 1022 -1743 1038
rect -1617 1072 -1551 1088
rect -1617 1038 -1601 1072
rect -1567 1038 -1551 1072
rect -1791 1000 -1761 1022
rect -1695 1000 -1665 1026
rect -1617 1022 -1551 1038
rect -1425 1072 -1359 1088
rect -1425 1038 -1409 1072
rect -1375 1038 -1359 1072
rect -1599 1000 -1569 1022
rect -1503 1000 -1473 1026
rect -1425 1022 -1359 1038
rect -1233 1072 -1167 1088
rect -1233 1038 -1217 1072
rect -1183 1038 -1167 1072
rect -1407 1000 -1377 1022
rect -1311 1000 -1281 1026
rect -1233 1022 -1167 1038
rect -1041 1072 -975 1088
rect -1041 1038 -1025 1072
rect -991 1038 -975 1072
rect -1215 1000 -1185 1022
rect -1119 1000 -1089 1026
rect -1041 1022 -975 1038
rect -849 1072 -783 1088
rect -849 1038 -833 1072
rect -799 1038 -783 1072
rect -1023 1000 -993 1022
rect -927 1000 -897 1026
rect -849 1022 -783 1038
rect -657 1072 -591 1088
rect -657 1038 -641 1072
rect -607 1038 -591 1072
rect -831 1000 -801 1022
rect -735 1000 -705 1026
rect -657 1022 -591 1038
rect -465 1072 -399 1088
rect -465 1038 -449 1072
rect -415 1038 -399 1072
rect -639 1000 -609 1022
rect -543 1000 -513 1026
rect -465 1022 -399 1038
rect -273 1072 -207 1088
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -447 1000 -417 1022
rect -351 1000 -321 1026
rect -273 1022 -207 1038
rect -81 1072 -15 1088
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect -255 1000 -225 1022
rect -159 1000 -129 1026
rect -81 1022 -15 1038
rect 111 1072 177 1088
rect 111 1038 127 1072
rect 161 1038 177 1072
rect -63 1000 -33 1022
rect 33 1000 63 1026
rect 111 1022 177 1038
rect 303 1072 369 1088
rect 303 1038 319 1072
rect 353 1038 369 1072
rect 129 1000 159 1022
rect 225 1000 255 1026
rect 303 1022 369 1038
rect 495 1072 561 1088
rect 495 1038 511 1072
rect 545 1038 561 1072
rect 321 1000 351 1022
rect 417 1000 447 1026
rect 495 1022 561 1038
rect 687 1072 753 1088
rect 687 1038 703 1072
rect 737 1038 753 1072
rect 513 1000 543 1022
rect 609 1000 639 1026
rect 687 1022 753 1038
rect 879 1072 945 1088
rect 879 1038 895 1072
rect 929 1038 945 1072
rect 705 1000 735 1022
rect 801 1000 831 1026
rect 879 1022 945 1038
rect 1071 1072 1137 1088
rect 1071 1038 1087 1072
rect 1121 1038 1137 1072
rect 897 1000 927 1022
rect 993 1000 1023 1026
rect 1071 1022 1137 1038
rect 1263 1072 1329 1088
rect 1263 1038 1279 1072
rect 1313 1038 1329 1072
rect 1089 1000 1119 1022
rect 1185 1000 1215 1026
rect 1263 1022 1329 1038
rect 1455 1072 1521 1088
rect 1455 1038 1471 1072
rect 1505 1038 1521 1072
rect 1281 1000 1311 1022
rect 1377 1000 1407 1026
rect 1455 1022 1521 1038
rect 1647 1072 1713 1088
rect 1647 1038 1663 1072
rect 1697 1038 1713 1072
rect 1473 1000 1503 1022
rect 1569 1000 1599 1026
rect 1647 1022 1713 1038
rect 1839 1072 1905 1088
rect 1839 1038 1855 1072
rect 1889 1038 1905 1072
rect 1665 1000 1695 1022
rect 1761 1000 1791 1026
rect 1839 1022 1905 1038
rect 2031 1072 2097 1088
rect 2031 1038 2047 1072
rect 2081 1038 2097 1072
rect 1857 1000 1887 1022
rect 1953 1000 1983 1026
rect 2031 1022 2097 1038
rect 2223 1072 2289 1088
rect 2223 1038 2239 1072
rect 2273 1038 2289 1072
rect 2049 1000 2079 1022
rect 2145 1000 2175 1026
rect 2223 1022 2289 1038
rect 2415 1072 2481 1088
rect 2415 1038 2431 1072
rect 2465 1038 2481 1072
rect 2241 1000 2271 1022
rect 2337 1000 2367 1026
rect 2415 1022 2481 1038
rect 2607 1072 2673 1088
rect 2607 1038 2623 1072
rect 2657 1038 2673 1072
rect 2433 1000 2463 1022
rect 2529 1000 2559 1026
rect 2607 1022 2673 1038
rect 2799 1072 2865 1088
rect 2799 1038 2815 1072
rect 2849 1038 2865 1072
rect 2625 1000 2655 1022
rect 2721 1000 2751 1026
rect 2799 1022 2865 1038
rect 2991 1072 3057 1088
rect 2991 1038 3007 1072
rect 3041 1038 3057 1072
rect 2817 1000 2847 1022
rect 2913 1000 2943 1026
rect 2991 1022 3057 1038
rect 3183 1072 3249 1088
rect 3183 1038 3199 1072
rect 3233 1038 3249 1072
rect 3009 1000 3039 1022
rect 3105 1000 3135 1026
rect 3183 1022 3249 1038
rect 3375 1072 3441 1088
rect 3375 1038 3391 1072
rect 3425 1038 3441 1072
rect 3201 1000 3231 1022
rect 3297 1000 3327 1026
rect 3375 1022 3441 1038
rect 3567 1072 3633 1088
rect 3567 1038 3583 1072
rect 3617 1038 3633 1072
rect 3393 1000 3423 1022
rect 3489 1000 3519 1026
rect 3567 1022 3633 1038
rect 3759 1072 3825 1088
rect 3759 1038 3775 1072
rect 3809 1038 3825 1072
rect 3585 1000 3615 1022
rect 3681 1000 3711 1026
rect 3759 1022 3825 1038
rect 3951 1072 4017 1088
rect 3951 1038 3967 1072
rect 4001 1038 4017 1072
rect 3777 1000 3807 1022
rect 3873 1000 3903 1026
rect 3951 1022 4017 1038
rect 4143 1072 4209 1088
rect 4143 1038 4159 1072
rect 4193 1038 4209 1072
rect 3969 1000 3999 1022
rect 4065 1000 4095 1026
rect 4143 1022 4209 1038
rect 4335 1072 4401 1088
rect 4335 1038 4351 1072
rect 4385 1038 4401 1072
rect 4161 1000 4191 1022
rect 4257 1000 4287 1026
rect 4335 1022 4401 1038
rect 4527 1072 4593 1088
rect 4527 1038 4543 1072
rect 4577 1038 4593 1072
rect 4353 1000 4383 1022
rect 4449 1000 4479 1026
rect 4527 1022 4593 1038
rect 4719 1072 4785 1088
rect 4719 1038 4735 1072
rect 4769 1038 4785 1072
rect 4545 1000 4575 1022
rect 4641 1000 4671 1026
rect 4719 1022 4785 1038
rect 4737 1000 4767 1022
rect -4767 -1022 -4737 -1000
rect -4785 -1038 -4719 -1022
rect -4671 -1026 -4641 -1000
rect -4575 -1022 -4545 -1000
rect -4785 -1072 -4769 -1038
rect -4735 -1072 -4719 -1038
rect -4785 -1088 -4719 -1072
rect -4593 -1038 -4527 -1022
rect -4479 -1026 -4449 -1000
rect -4383 -1022 -4353 -1000
rect -4593 -1072 -4577 -1038
rect -4543 -1072 -4527 -1038
rect -4593 -1088 -4527 -1072
rect -4401 -1038 -4335 -1022
rect -4287 -1026 -4257 -1000
rect -4191 -1022 -4161 -1000
rect -4401 -1072 -4385 -1038
rect -4351 -1072 -4335 -1038
rect -4401 -1088 -4335 -1072
rect -4209 -1038 -4143 -1022
rect -4095 -1026 -4065 -1000
rect -3999 -1022 -3969 -1000
rect -4209 -1072 -4193 -1038
rect -4159 -1072 -4143 -1038
rect -4209 -1088 -4143 -1072
rect -4017 -1038 -3951 -1022
rect -3903 -1026 -3873 -1000
rect -3807 -1022 -3777 -1000
rect -4017 -1072 -4001 -1038
rect -3967 -1072 -3951 -1038
rect -4017 -1088 -3951 -1072
rect -3825 -1038 -3759 -1022
rect -3711 -1026 -3681 -1000
rect -3615 -1022 -3585 -1000
rect -3825 -1072 -3809 -1038
rect -3775 -1072 -3759 -1038
rect -3825 -1088 -3759 -1072
rect -3633 -1038 -3567 -1022
rect -3519 -1026 -3489 -1000
rect -3423 -1022 -3393 -1000
rect -3633 -1072 -3617 -1038
rect -3583 -1072 -3567 -1038
rect -3633 -1088 -3567 -1072
rect -3441 -1038 -3375 -1022
rect -3327 -1026 -3297 -1000
rect -3231 -1022 -3201 -1000
rect -3441 -1072 -3425 -1038
rect -3391 -1072 -3375 -1038
rect -3441 -1088 -3375 -1072
rect -3249 -1038 -3183 -1022
rect -3135 -1026 -3105 -1000
rect -3039 -1022 -3009 -1000
rect -3249 -1072 -3233 -1038
rect -3199 -1072 -3183 -1038
rect -3249 -1088 -3183 -1072
rect -3057 -1038 -2991 -1022
rect -2943 -1026 -2913 -1000
rect -2847 -1022 -2817 -1000
rect -3057 -1072 -3041 -1038
rect -3007 -1072 -2991 -1038
rect -3057 -1088 -2991 -1072
rect -2865 -1038 -2799 -1022
rect -2751 -1026 -2721 -1000
rect -2655 -1022 -2625 -1000
rect -2865 -1072 -2849 -1038
rect -2815 -1072 -2799 -1038
rect -2865 -1088 -2799 -1072
rect -2673 -1038 -2607 -1022
rect -2559 -1026 -2529 -1000
rect -2463 -1022 -2433 -1000
rect -2673 -1072 -2657 -1038
rect -2623 -1072 -2607 -1038
rect -2673 -1088 -2607 -1072
rect -2481 -1038 -2415 -1022
rect -2367 -1026 -2337 -1000
rect -2271 -1022 -2241 -1000
rect -2481 -1072 -2465 -1038
rect -2431 -1072 -2415 -1038
rect -2481 -1088 -2415 -1072
rect -2289 -1038 -2223 -1022
rect -2175 -1026 -2145 -1000
rect -2079 -1022 -2049 -1000
rect -2289 -1072 -2273 -1038
rect -2239 -1072 -2223 -1038
rect -2289 -1088 -2223 -1072
rect -2097 -1038 -2031 -1022
rect -1983 -1026 -1953 -1000
rect -1887 -1022 -1857 -1000
rect -2097 -1072 -2081 -1038
rect -2047 -1072 -2031 -1038
rect -2097 -1088 -2031 -1072
rect -1905 -1038 -1839 -1022
rect -1791 -1026 -1761 -1000
rect -1695 -1022 -1665 -1000
rect -1905 -1072 -1889 -1038
rect -1855 -1072 -1839 -1038
rect -1905 -1088 -1839 -1072
rect -1713 -1038 -1647 -1022
rect -1599 -1026 -1569 -1000
rect -1503 -1022 -1473 -1000
rect -1713 -1072 -1697 -1038
rect -1663 -1072 -1647 -1038
rect -1713 -1088 -1647 -1072
rect -1521 -1038 -1455 -1022
rect -1407 -1026 -1377 -1000
rect -1311 -1022 -1281 -1000
rect -1521 -1072 -1505 -1038
rect -1471 -1072 -1455 -1038
rect -1521 -1088 -1455 -1072
rect -1329 -1038 -1263 -1022
rect -1215 -1026 -1185 -1000
rect -1119 -1022 -1089 -1000
rect -1329 -1072 -1313 -1038
rect -1279 -1072 -1263 -1038
rect -1329 -1088 -1263 -1072
rect -1137 -1038 -1071 -1022
rect -1023 -1026 -993 -1000
rect -927 -1022 -897 -1000
rect -1137 -1072 -1121 -1038
rect -1087 -1072 -1071 -1038
rect -1137 -1088 -1071 -1072
rect -945 -1038 -879 -1022
rect -831 -1026 -801 -1000
rect -735 -1022 -705 -1000
rect -945 -1072 -929 -1038
rect -895 -1072 -879 -1038
rect -945 -1088 -879 -1072
rect -753 -1038 -687 -1022
rect -639 -1026 -609 -1000
rect -543 -1022 -513 -1000
rect -753 -1072 -737 -1038
rect -703 -1072 -687 -1038
rect -753 -1088 -687 -1072
rect -561 -1038 -495 -1022
rect -447 -1026 -417 -1000
rect -351 -1022 -321 -1000
rect -561 -1072 -545 -1038
rect -511 -1072 -495 -1038
rect -561 -1088 -495 -1072
rect -369 -1038 -303 -1022
rect -255 -1026 -225 -1000
rect -159 -1022 -129 -1000
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -369 -1088 -303 -1072
rect -177 -1038 -111 -1022
rect -63 -1026 -33 -1000
rect 33 -1022 63 -1000
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect -177 -1088 -111 -1072
rect 15 -1038 81 -1022
rect 129 -1026 159 -1000
rect 225 -1022 255 -1000
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 15 -1088 81 -1072
rect 207 -1038 273 -1022
rect 321 -1026 351 -1000
rect 417 -1022 447 -1000
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 207 -1088 273 -1072
rect 399 -1038 465 -1022
rect 513 -1026 543 -1000
rect 609 -1022 639 -1000
rect 399 -1072 415 -1038
rect 449 -1072 465 -1038
rect 399 -1088 465 -1072
rect 591 -1038 657 -1022
rect 705 -1026 735 -1000
rect 801 -1022 831 -1000
rect 591 -1072 607 -1038
rect 641 -1072 657 -1038
rect 591 -1088 657 -1072
rect 783 -1038 849 -1022
rect 897 -1026 927 -1000
rect 993 -1022 1023 -1000
rect 783 -1072 799 -1038
rect 833 -1072 849 -1038
rect 783 -1088 849 -1072
rect 975 -1038 1041 -1022
rect 1089 -1026 1119 -1000
rect 1185 -1022 1215 -1000
rect 975 -1072 991 -1038
rect 1025 -1072 1041 -1038
rect 975 -1088 1041 -1072
rect 1167 -1038 1233 -1022
rect 1281 -1026 1311 -1000
rect 1377 -1022 1407 -1000
rect 1167 -1072 1183 -1038
rect 1217 -1072 1233 -1038
rect 1167 -1088 1233 -1072
rect 1359 -1038 1425 -1022
rect 1473 -1026 1503 -1000
rect 1569 -1022 1599 -1000
rect 1359 -1072 1375 -1038
rect 1409 -1072 1425 -1038
rect 1359 -1088 1425 -1072
rect 1551 -1038 1617 -1022
rect 1665 -1026 1695 -1000
rect 1761 -1022 1791 -1000
rect 1551 -1072 1567 -1038
rect 1601 -1072 1617 -1038
rect 1551 -1088 1617 -1072
rect 1743 -1038 1809 -1022
rect 1857 -1026 1887 -1000
rect 1953 -1022 1983 -1000
rect 1743 -1072 1759 -1038
rect 1793 -1072 1809 -1038
rect 1743 -1088 1809 -1072
rect 1935 -1038 2001 -1022
rect 2049 -1026 2079 -1000
rect 2145 -1022 2175 -1000
rect 1935 -1072 1951 -1038
rect 1985 -1072 2001 -1038
rect 1935 -1088 2001 -1072
rect 2127 -1038 2193 -1022
rect 2241 -1026 2271 -1000
rect 2337 -1022 2367 -1000
rect 2127 -1072 2143 -1038
rect 2177 -1072 2193 -1038
rect 2127 -1088 2193 -1072
rect 2319 -1038 2385 -1022
rect 2433 -1026 2463 -1000
rect 2529 -1022 2559 -1000
rect 2319 -1072 2335 -1038
rect 2369 -1072 2385 -1038
rect 2319 -1088 2385 -1072
rect 2511 -1038 2577 -1022
rect 2625 -1026 2655 -1000
rect 2721 -1022 2751 -1000
rect 2511 -1072 2527 -1038
rect 2561 -1072 2577 -1038
rect 2511 -1088 2577 -1072
rect 2703 -1038 2769 -1022
rect 2817 -1026 2847 -1000
rect 2913 -1022 2943 -1000
rect 2703 -1072 2719 -1038
rect 2753 -1072 2769 -1038
rect 2703 -1088 2769 -1072
rect 2895 -1038 2961 -1022
rect 3009 -1026 3039 -1000
rect 3105 -1022 3135 -1000
rect 2895 -1072 2911 -1038
rect 2945 -1072 2961 -1038
rect 2895 -1088 2961 -1072
rect 3087 -1038 3153 -1022
rect 3201 -1026 3231 -1000
rect 3297 -1022 3327 -1000
rect 3087 -1072 3103 -1038
rect 3137 -1072 3153 -1038
rect 3087 -1088 3153 -1072
rect 3279 -1038 3345 -1022
rect 3393 -1026 3423 -1000
rect 3489 -1022 3519 -1000
rect 3279 -1072 3295 -1038
rect 3329 -1072 3345 -1038
rect 3279 -1088 3345 -1072
rect 3471 -1038 3537 -1022
rect 3585 -1026 3615 -1000
rect 3681 -1022 3711 -1000
rect 3471 -1072 3487 -1038
rect 3521 -1072 3537 -1038
rect 3471 -1088 3537 -1072
rect 3663 -1038 3729 -1022
rect 3777 -1026 3807 -1000
rect 3873 -1022 3903 -1000
rect 3663 -1072 3679 -1038
rect 3713 -1072 3729 -1038
rect 3663 -1088 3729 -1072
rect 3855 -1038 3921 -1022
rect 3969 -1026 3999 -1000
rect 4065 -1022 4095 -1000
rect 3855 -1072 3871 -1038
rect 3905 -1072 3921 -1038
rect 3855 -1088 3921 -1072
rect 4047 -1038 4113 -1022
rect 4161 -1026 4191 -1000
rect 4257 -1022 4287 -1000
rect 4047 -1072 4063 -1038
rect 4097 -1072 4113 -1038
rect 4047 -1088 4113 -1072
rect 4239 -1038 4305 -1022
rect 4353 -1026 4383 -1000
rect 4449 -1022 4479 -1000
rect 4239 -1072 4255 -1038
rect 4289 -1072 4305 -1038
rect 4239 -1088 4305 -1072
rect 4431 -1038 4497 -1022
rect 4545 -1026 4575 -1000
rect 4641 -1022 4671 -1000
rect 4431 -1072 4447 -1038
rect 4481 -1072 4497 -1038
rect 4431 -1088 4497 -1072
rect 4623 -1038 4689 -1022
rect 4737 -1026 4767 -1000
rect 4623 -1072 4639 -1038
rect 4673 -1072 4689 -1038
rect 4623 -1088 4689 -1072
<< polycont >>
rect -4673 1038 -4639 1072
rect -4481 1038 -4447 1072
rect -4289 1038 -4255 1072
rect -4097 1038 -4063 1072
rect -3905 1038 -3871 1072
rect -3713 1038 -3679 1072
rect -3521 1038 -3487 1072
rect -3329 1038 -3295 1072
rect -3137 1038 -3103 1072
rect -2945 1038 -2911 1072
rect -2753 1038 -2719 1072
rect -2561 1038 -2527 1072
rect -2369 1038 -2335 1072
rect -2177 1038 -2143 1072
rect -1985 1038 -1951 1072
rect -1793 1038 -1759 1072
rect -1601 1038 -1567 1072
rect -1409 1038 -1375 1072
rect -1217 1038 -1183 1072
rect -1025 1038 -991 1072
rect -833 1038 -799 1072
rect -641 1038 -607 1072
rect -449 1038 -415 1072
rect -257 1038 -223 1072
rect -65 1038 -31 1072
rect 127 1038 161 1072
rect 319 1038 353 1072
rect 511 1038 545 1072
rect 703 1038 737 1072
rect 895 1038 929 1072
rect 1087 1038 1121 1072
rect 1279 1038 1313 1072
rect 1471 1038 1505 1072
rect 1663 1038 1697 1072
rect 1855 1038 1889 1072
rect 2047 1038 2081 1072
rect 2239 1038 2273 1072
rect 2431 1038 2465 1072
rect 2623 1038 2657 1072
rect 2815 1038 2849 1072
rect 3007 1038 3041 1072
rect 3199 1038 3233 1072
rect 3391 1038 3425 1072
rect 3583 1038 3617 1072
rect 3775 1038 3809 1072
rect 3967 1038 4001 1072
rect 4159 1038 4193 1072
rect 4351 1038 4385 1072
rect 4543 1038 4577 1072
rect 4735 1038 4769 1072
rect -4769 -1072 -4735 -1038
rect -4577 -1072 -4543 -1038
rect -4385 -1072 -4351 -1038
rect -4193 -1072 -4159 -1038
rect -4001 -1072 -3967 -1038
rect -3809 -1072 -3775 -1038
rect -3617 -1072 -3583 -1038
rect -3425 -1072 -3391 -1038
rect -3233 -1072 -3199 -1038
rect -3041 -1072 -3007 -1038
rect -2849 -1072 -2815 -1038
rect -2657 -1072 -2623 -1038
rect -2465 -1072 -2431 -1038
rect -2273 -1072 -2239 -1038
rect -2081 -1072 -2047 -1038
rect -1889 -1072 -1855 -1038
rect -1697 -1072 -1663 -1038
rect -1505 -1072 -1471 -1038
rect -1313 -1072 -1279 -1038
rect -1121 -1072 -1087 -1038
rect -929 -1072 -895 -1038
rect -737 -1072 -703 -1038
rect -545 -1072 -511 -1038
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
rect 415 -1072 449 -1038
rect 607 -1072 641 -1038
rect 799 -1072 833 -1038
rect 991 -1072 1025 -1038
rect 1183 -1072 1217 -1038
rect 1375 -1072 1409 -1038
rect 1567 -1072 1601 -1038
rect 1759 -1072 1793 -1038
rect 1951 -1072 1985 -1038
rect 2143 -1072 2177 -1038
rect 2335 -1072 2369 -1038
rect 2527 -1072 2561 -1038
rect 2719 -1072 2753 -1038
rect 2911 -1072 2945 -1038
rect 3103 -1072 3137 -1038
rect 3295 -1072 3329 -1038
rect 3487 -1072 3521 -1038
rect 3679 -1072 3713 -1038
rect 3871 -1072 3905 -1038
rect 4063 -1072 4097 -1038
rect 4255 -1072 4289 -1038
rect 4447 -1072 4481 -1038
rect 4639 -1072 4673 -1038
<< locali >>
rect -4931 1140 -4835 1174
rect 4835 1140 4931 1174
rect -4931 1078 -4897 1140
rect 4897 1078 4931 1140
rect -4689 1038 -4673 1072
rect -4639 1038 -4623 1072
rect -4497 1038 -4481 1072
rect -4447 1038 -4431 1072
rect -4305 1038 -4289 1072
rect -4255 1038 -4239 1072
rect -4113 1038 -4097 1072
rect -4063 1038 -4047 1072
rect -3921 1038 -3905 1072
rect -3871 1038 -3855 1072
rect -3729 1038 -3713 1072
rect -3679 1038 -3663 1072
rect -3537 1038 -3521 1072
rect -3487 1038 -3471 1072
rect -3345 1038 -3329 1072
rect -3295 1038 -3279 1072
rect -3153 1038 -3137 1072
rect -3103 1038 -3087 1072
rect -2961 1038 -2945 1072
rect -2911 1038 -2895 1072
rect -2769 1038 -2753 1072
rect -2719 1038 -2703 1072
rect -2577 1038 -2561 1072
rect -2527 1038 -2511 1072
rect -2385 1038 -2369 1072
rect -2335 1038 -2319 1072
rect -2193 1038 -2177 1072
rect -2143 1038 -2127 1072
rect -2001 1038 -1985 1072
rect -1951 1038 -1935 1072
rect -1809 1038 -1793 1072
rect -1759 1038 -1743 1072
rect -1617 1038 -1601 1072
rect -1567 1038 -1551 1072
rect -1425 1038 -1409 1072
rect -1375 1038 -1359 1072
rect -1233 1038 -1217 1072
rect -1183 1038 -1167 1072
rect -1041 1038 -1025 1072
rect -991 1038 -975 1072
rect -849 1038 -833 1072
rect -799 1038 -783 1072
rect -657 1038 -641 1072
rect -607 1038 -591 1072
rect -465 1038 -449 1072
rect -415 1038 -399 1072
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect 111 1038 127 1072
rect 161 1038 177 1072
rect 303 1038 319 1072
rect 353 1038 369 1072
rect 495 1038 511 1072
rect 545 1038 561 1072
rect 687 1038 703 1072
rect 737 1038 753 1072
rect 879 1038 895 1072
rect 929 1038 945 1072
rect 1071 1038 1087 1072
rect 1121 1038 1137 1072
rect 1263 1038 1279 1072
rect 1313 1038 1329 1072
rect 1455 1038 1471 1072
rect 1505 1038 1521 1072
rect 1647 1038 1663 1072
rect 1697 1038 1713 1072
rect 1839 1038 1855 1072
rect 1889 1038 1905 1072
rect 2031 1038 2047 1072
rect 2081 1038 2097 1072
rect 2223 1038 2239 1072
rect 2273 1038 2289 1072
rect 2415 1038 2431 1072
rect 2465 1038 2481 1072
rect 2607 1038 2623 1072
rect 2657 1038 2673 1072
rect 2799 1038 2815 1072
rect 2849 1038 2865 1072
rect 2991 1038 3007 1072
rect 3041 1038 3057 1072
rect 3183 1038 3199 1072
rect 3233 1038 3249 1072
rect 3375 1038 3391 1072
rect 3425 1038 3441 1072
rect 3567 1038 3583 1072
rect 3617 1038 3633 1072
rect 3759 1038 3775 1072
rect 3809 1038 3825 1072
rect 3951 1038 3967 1072
rect 4001 1038 4017 1072
rect 4143 1038 4159 1072
rect 4193 1038 4209 1072
rect 4335 1038 4351 1072
rect 4385 1038 4401 1072
rect 4527 1038 4543 1072
rect 4577 1038 4593 1072
rect 4719 1038 4735 1072
rect 4769 1038 4785 1072
rect -4817 988 -4783 1004
rect -4817 -1004 -4783 -988
rect -4721 988 -4687 1004
rect -4721 -1004 -4687 -988
rect -4625 988 -4591 1004
rect -4625 -1004 -4591 -988
rect -4529 988 -4495 1004
rect -4529 -1004 -4495 -988
rect -4433 988 -4399 1004
rect -4433 -1004 -4399 -988
rect -4337 988 -4303 1004
rect -4337 -1004 -4303 -988
rect -4241 988 -4207 1004
rect -4241 -1004 -4207 -988
rect -4145 988 -4111 1004
rect -4145 -1004 -4111 -988
rect -4049 988 -4015 1004
rect -4049 -1004 -4015 -988
rect -3953 988 -3919 1004
rect -3953 -1004 -3919 -988
rect -3857 988 -3823 1004
rect -3857 -1004 -3823 -988
rect -3761 988 -3727 1004
rect -3761 -1004 -3727 -988
rect -3665 988 -3631 1004
rect -3665 -1004 -3631 -988
rect -3569 988 -3535 1004
rect -3569 -1004 -3535 -988
rect -3473 988 -3439 1004
rect -3473 -1004 -3439 -988
rect -3377 988 -3343 1004
rect -3377 -1004 -3343 -988
rect -3281 988 -3247 1004
rect -3281 -1004 -3247 -988
rect -3185 988 -3151 1004
rect -3185 -1004 -3151 -988
rect -3089 988 -3055 1004
rect -3089 -1004 -3055 -988
rect -2993 988 -2959 1004
rect -2993 -1004 -2959 -988
rect -2897 988 -2863 1004
rect -2897 -1004 -2863 -988
rect -2801 988 -2767 1004
rect -2801 -1004 -2767 -988
rect -2705 988 -2671 1004
rect -2705 -1004 -2671 -988
rect -2609 988 -2575 1004
rect -2609 -1004 -2575 -988
rect -2513 988 -2479 1004
rect -2513 -1004 -2479 -988
rect -2417 988 -2383 1004
rect -2417 -1004 -2383 -988
rect -2321 988 -2287 1004
rect -2321 -1004 -2287 -988
rect -2225 988 -2191 1004
rect -2225 -1004 -2191 -988
rect -2129 988 -2095 1004
rect -2129 -1004 -2095 -988
rect -2033 988 -1999 1004
rect -2033 -1004 -1999 -988
rect -1937 988 -1903 1004
rect -1937 -1004 -1903 -988
rect -1841 988 -1807 1004
rect -1841 -1004 -1807 -988
rect -1745 988 -1711 1004
rect -1745 -1004 -1711 -988
rect -1649 988 -1615 1004
rect -1649 -1004 -1615 -988
rect -1553 988 -1519 1004
rect -1553 -1004 -1519 -988
rect -1457 988 -1423 1004
rect -1457 -1004 -1423 -988
rect -1361 988 -1327 1004
rect -1361 -1004 -1327 -988
rect -1265 988 -1231 1004
rect -1265 -1004 -1231 -988
rect -1169 988 -1135 1004
rect -1169 -1004 -1135 -988
rect -1073 988 -1039 1004
rect -1073 -1004 -1039 -988
rect -977 988 -943 1004
rect -977 -1004 -943 -988
rect -881 988 -847 1004
rect -881 -1004 -847 -988
rect -785 988 -751 1004
rect -785 -1004 -751 -988
rect -689 988 -655 1004
rect -689 -1004 -655 -988
rect -593 988 -559 1004
rect -593 -1004 -559 -988
rect -497 988 -463 1004
rect -497 -1004 -463 -988
rect -401 988 -367 1004
rect -401 -1004 -367 -988
rect -305 988 -271 1004
rect -305 -1004 -271 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 271 988 305 1004
rect 271 -1004 305 -988
rect 367 988 401 1004
rect 367 -1004 401 -988
rect 463 988 497 1004
rect 463 -1004 497 -988
rect 559 988 593 1004
rect 559 -1004 593 -988
rect 655 988 689 1004
rect 655 -1004 689 -988
rect 751 988 785 1004
rect 751 -1004 785 -988
rect 847 988 881 1004
rect 847 -1004 881 -988
rect 943 988 977 1004
rect 943 -1004 977 -988
rect 1039 988 1073 1004
rect 1039 -1004 1073 -988
rect 1135 988 1169 1004
rect 1135 -1004 1169 -988
rect 1231 988 1265 1004
rect 1231 -1004 1265 -988
rect 1327 988 1361 1004
rect 1327 -1004 1361 -988
rect 1423 988 1457 1004
rect 1423 -1004 1457 -988
rect 1519 988 1553 1004
rect 1519 -1004 1553 -988
rect 1615 988 1649 1004
rect 1615 -1004 1649 -988
rect 1711 988 1745 1004
rect 1711 -1004 1745 -988
rect 1807 988 1841 1004
rect 1807 -1004 1841 -988
rect 1903 988 1937 1004
rect 1903 -1004 1937 -988
rect 1999 988 2033 1004
rect 1999 -1004 2033 -988
rect 2095 988 2129 1004
rect 2095 -1004 2129 -988
rect 2191 988 2225 1004
rect 2191 -1004 2225 -988
rect 2287 988 2321 1004
rect 2287 -1004 2321 -988
rect 2383 988 2417 1004
rect 2383 -1004 2417 -988
rect 2479 988 2513 1004
rect 2479 -1004 2513 -988
rect 2575 988 2609 1004
rect 2575 -1004 2609 -988
rect 2671 988 2705 1004
rect 2671 -1004 2705 -988
rect 2767 988 2801 1004
rect 2767 -1004 2801 -988
rect 2863 988 2897 1004
rect 2863 -1004 2897 -988
rect 2959 988 2993 1004
rect 2959 -1004 2993 -988
rect 3055 988 3089 1004
rect 3055 -1004 3089 -988
rect 3151 988 3185 1004
rect 3151 -1004 3185 -988
rect 3247 988 3281 1004
rect 3247 -1004 3281 -988
rect 3343 988 3377 1004
rect 3343 -1004 3377 -988
rect 3439 988 3473 1004
rect 3439 -1004 3473 -988
rect 3535 988 3569 1004
rect 3535 -1004 3569 -988
rect 3631 988 3665 1004
rect 3631 -1004 3665 -988
rect 3727 988 3761 1004
rect 3727 -1004 3761 -988
rect 3823 988 3857 1004
rect 3823 -1004 3857 -988
rect 3919 988 3953 1004
rect 3919 -1004 3953 -988
rect 4015 988 4049 1004
rect 4015 -1004 4049 -988
rect 4111 988 4145 1004
rect 4111 -1004 4145 -988
rect 4207 988 4241 1004
rect 4207 -1004 4241 -988
rect 4303 988 4337 1004
rect 4303 -1004 4337 -988
rect 4399 988 4433 1004
rect 4399 -1004 4433 -988
rect 4495 988 4529 1004
rect 4495 -1004 4529 -988
rect 4591 988 4625 1004
rect 4591 -1004 4625 -988
rect 4687 988 4721 1004
rect 4687 -1004 4721 -988
rect 4783 988 4817 1004
rect 4783 -1004 4817 -988
rect -4785 -1072 -4769 -1038
rect -4735 -1072 -4719 -1038
rect -4593 -1072 -4577 -1038
rect -4543 -1072 -4527 -1038
rect -4401 -1072 -4385 -1038
rect -4351 -1072 -4335 -1038
rect -4209 -1072 -4193 -1038
rect -4159 -1072 -4143 -1038
rect -4017 -1072 -4001 -1038
rect -3967 -1072 -3951 -1038
rect -3825 -1072 -3809 -1038
rect -3775 -1072 -3759 -1038
rect -3633 -1072 -3617 -1038
rect -3583 -1072 -3567 -1038
rect -3441 -1072 -3425 -1038
rect -3391 -1072 -3375 -1038
rect -3249 -1072 -3233 -1038
rect -3199 -1072 -3183 -1038
rect -3057 -1072 -3041 -1038
rect -3007 -1072 -2991 -1038
rect -2865 -1072 -2849 -1038
rect -2815 -1072 -2799 -1038
rect -2673 -1072 -2657 -1038
rect -2623 -1072 -2607 -1038
rect -2481 -1072 -2465 -1038
rect -2431 -1072 -2415 -1038
rect -2289 -1072 -2273 -1038
rect -2239 -1072 -2223 -1038
rect -2097 -1072 -2081 -1038
rect -2047 -1072 -2031 -1038
rect -1905 -1072 -1889 -1038
rect -1855 -1072 -1839 -1038
rect -1713 -1072 -1697 -1038
rect -1663 -1072 -1647 -1038
rect -1521 -1072 -1505 -1038
rect -1471 -1072 -1455 -1038
rect -1329 -1072 -1313 -1038
rect -1279 -1072 -1263 -1038
rect -1137 -1072 -1121 -1038
rect -1087 -1072 -1071 -1038
rect -945 -1072 -929 -1038
rect -895 -1072 -879 -1038
rect -753 -1072 -737 -1038
rect -703 -1072 -687 -1038
rect -561 -1072 -545 -1038
rect -511 -1072 -495 -1038
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 399 -1072 415 -1038
rect 449 -1072 465 -1038
rect 591 -1072 607 -1038
rect 641 -1072 657 -1038
rect 783 -1072 799 -1038
rect 833 -1072 849 -1038
rect 975 -1072 991 -1038
rect 1025 -1072 1041 -1038
rect 1167 -1072 1183 -1038
rect 1217 -1072 1233 -1038
rect 1359 -1072 1375 -1038
rect 1409 -1072 1425 -1038
rect 1551 -1072 1567 -1038
rect 1601 -1072 1617 -1038
rect 1743 -1072 1759 -1038
rect 1793 -1072 1809 -1038
rect 1935 -1072 1951 -1038
rect 1985 -1072 2001 -1038
rect 2127 -1072 2143 -1038
rect 2177 -1072 2193 -1038
rect 2319 -1072 2335 -1038
rect 2369 -1072 2385 -1038
rect 2511 -1072 2527 -1038
rect 2561 -1072 2577 -1038
rect 2703 -1072 2719 -1038
rect 2753 -1072 2769 -1038
rect 2895 -1072 2911 -1038
rect 2945 -1072 2961 -1038
rect 3087 -1072 3103 -1038
rect 3137 -1072 3153 -1038
rect 3279 -1072 3295 -1038
rect 3329 -1072 3345 -1038
rect 3471 -1072 3487 -1038
rect 3521 -1072 3537 -1038
rect 3663 -1072 3679 -1038
rect 3713 -1072 3729 -1038
rect 3855 -1072 3871 -1038
rect 3905 -1072 3921 -1038
rect 4047 -1072 4063 -1038
rect 4097 -1072 4113 -1038
rect 4239 -1072 4255 -1038
rect 4289 -1072 4305 -1038
rect 4431 -1072 4447 -1038
rect 4481 -1072 4497 -1038
rect 4623 -1072 4639 -1038
rect 4673 -1072 4689 -1038
rect -4931 -1140 -4897 -1078
rect 4897 -1140 4931 -1078
rect -4931 -1174 -4835 -1140
rect 4835 -1174 4931 -1140
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -4914 -1157 4914 1157
string parameters w 10 l 0.150 m 1 nf 100 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
