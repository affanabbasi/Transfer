magic
tech sky130A
magscale 1 2
timestamp 1606578544
<< pwell >>
rect -201 -1057 201 1057
<< psubdiff >>
rect -165 987 -69 1021
rect 69 987 165 1021
rect -165 925 -131 987
rect 131 925 165 987
rect -165 -987 -131 -925
rect 131 -987 165 -925
rect -165 -1021 -69 -987
rect 69 -1021 165 -987
<< psubdiffcont >>
rect -69 987 69 1021
rect -165 -925 -131 925
rect 131 -925 165 925
rect -69 -1021 69 -987
<< xpolycontact >>
rect -35 459 35 891
rect -35 -891 35 -459
<< ppolyres >>
rect -35 -459 35 459
<< locali >>
rect -165 987 -69 1021
rect 69 987 165 1021
rect -165 925 -131 987
rect 131 925 165 987
rect -165 -987 -131 -925
rect 131 -987 165 -925
rect -165 -1021 -69 -987
rect 69 -1021 165 -987
<< res0p35 >>
rect -37 -461 37 461
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string FIXED_BBOX -148 -1004 148 1004
string parameters w 0.350 l 4.59 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 4.303k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350
string library sky130
<< end >>
