magic
tech sky130A
magscale 1 2
timestamp 1606670916
<< nwell >>
rect -348 312 118 652
<< pwell >>
rect 430 -804 1100 -68
rect -1212 -1620 -468 -1576
rect 430 -1620 1100 -962
rect 1660 -1620 2404 -1476
rect -1212 -1638 2404 -1620
rect -1212 -1852 2404 -1796
rect -1212 -1952 1760 -1852
rect -504 -2936 1760 -1952
<< viali >>
rect 88 324 130 358
rect 226 324 268 358
rect 402 324 444 358
rect 764 324 806 358
rect 878 324 920 358
rect 1008 324 1050 358
rect -558 278 -522 312
rect -460 220 -426 254
rect 164 209 340 243
rect 801 210 977 244
rect 71 165 105 199
rect 399 165 433 199
rect 708 166 742 200
rect 238 120 272 156
rect 902 122 938 158
rect -1042 -670 -972 -238
rect -724 -670 -654 -238
rect -406 -670 -336 -238
rect -88 -670 -18 -238
rect 230 -670 300 -238
rect 884 -666 954 -234
rect 1202 -666 1272 -234
rect 1520 -666 1590 -234
rect 1838 -666 1908 -234
rect 2156 -666 2226 -234
rect -1042 -1502 -972 -1070
rect -724 -1502 -654 -1070
rect -406 -1502 -336 -1070
rect -88 -1502 -18 -1070
rect 230 -1502 300 -1070
rect 884 -1498 954 -1066
rect 1202 -1498 1272 -1066
rect 1520 -1498 1590 -1066
rect 1838 -1498 1908 -1066
rect 2156 -1498 2226 -1066
rect -720 -1638 -662 -1596
rect 1838 -1630 1896 -1588
rect 1836 -1848 1894 -1806
rect -724 -1900 -666 -1858
rect -1030 -2426 -960 -1994
rect -712 -2426 -642 -1994
rect 1834 -2372 1904 -1940
rect 2152 -2372 2222 -1940
rect 1336 -2596 1442 -2562
rect -232 -2638 -126 -2604
rect 1248 -2640 1282 -2606
rect -72 -2682 -38 -2648
rect 1336 -2684 1442 -2650
rect -232 -2726 -126 -2692
rect -548 -2806 -512 -2770
rect 1246 -2800 1304 -2764
rect 1370 -2800 1428 -2764
rect 1474 -2800 1532 -2764
rect -322 -2840 -264 -2804
rect -206 -2842 -148 -2806
rect -94 -2840 -36 -2804
rect 1702 -2824 1738 -2788
rect -546 -2896 -510 -2860
rect 1702 -2898 1738 -2862
rect -1030 -5058 -960 -4626
rect -712 -5058 -642 -4626
rect 1834 -5004 1904 -4572
rect 2152 -5004 2222 -4572
<< metal1 >>
rect 272 706 734 842
rect 272 648 411 706
rect -382 552 411 648
rect -130 534 411 552
rect 604 648 734 706
rect 604 534 1228 648
rect -130 358 1228 534
rect -1316 324 -1230 332
rect -1316 272 -1294 324
rect -1240 320 -1230 324
rect -130 324 88 358
rect 130 324 226 358
rect 268 324 402 358
rect 444 324 764 358
rect 806 324 878 358
rect 920 324 1008 358
rect 1050 324 1228 358
rect -1240 312 -502 320
rect -1240 278 -558 312
rect -522 278 -502 312
rect -130 300 1228 324
rect -1240 272 -502 278
rect -1316 256 -502 272
rect -472 254 -80 266
rect -472 220 -460 254
rect -426 220 -80 254
rect -472 216 -80 220
rect 150 243 356 300
rect -472 206 120 216
rect -130 199 120 206
rect 150 209 164 243
rect 340 209 356 243
rect 788 244 992 300
rect 150 200 356 209
rect 386 200 758 216
rect -130 165 71 199
rect 105 165 120 199
rect 386 199 708 200
rect -130 142 120 165
rect 214 156 310 166
rect 214 120 238 156
rect 272 120 310 156
rect 386 165 399 199
rect 433 166 708 199
rect 742 166 758 200
rect 788 210 801 244
rect 977 210 992 244
rect 788 198 992 210
rect 433 165 758 166
rect 386 150 758 165
rect 862 158 968 168
rect -1070 -238 -624 -220
rect -1070 -670 -1042 -238
rect -972 -670 -724 -238
rect -654 -670 -624 -238
rect -1070 -682 -624 -670
rect -442 -238 8 -206
rect -442 -670 -406 -238
rect -336 -670 -88 -238
rect -18 -670 8 -238
rect -442 -678 8 -670
rect 214 -238 310 120
rect 214 -670 230 -238
rect 300 -670 310 -238
rect 214 -684 310 -670
rect 862 122 902 158
rect 938 122 968 158
rect 862 -234 968 122
rect 862 -666 884 -234
rect 954 -666 968 -234
rect 862 -676 968 -666
rect 1184 -234 1614 -198
rect 1184 -666 1202 -234
rect 1272 -666 1520 -234
rect 1590 -666 1614 -234
rect 1184 -678 1614 -666
rect 1818 -234 2244 -224
rect 1818 -666 1838 -234
rect 1908 -666 2156 -234
rect 2226 -666 2244 -234
rect 1818 -680 2244 -666
rect -1064 -1070 -940 -1042
rect -1064 -1502 -1042 -1070
rect -972 -1502 -940 -1070
rect -1064 -1676 -940 -1502
rect -766 -1070 -302 -1042
rect -766 -1502 -724 -1070
rect -654 -1502 -406 -1070
rect -336 -1502 -302 -1070
rect -766 -1522 -302 -1502
rect -112 -1070 330 -1050
rect -112 -1502 -88 -1070
rect -18 -1502 230 -1070
rect 300 -1502 330 -1070
rect -112 -1528 330 -1502
rect 868 -1066 1298 -1046
rect 868 -1498 884 -1066
rect 954 -1498 1202 -1066
rect 1272 -1498 1298 -1066
rect 868 -1526 1298 -1498
rect 1504 -1066 1934 -1030
rect 1504 -1498 1520 -1066
rect 1590 -1498 1838 -1066
rect 1908 -1498 1934 -1066
rect 1504 -1510 1934 -1498
rect 2128 -1066 2256 -1038
rect 2128 -1498 2156 -1066
rect 2226 -1498 2256 -1066
rect -1090 -1696 -940 -1676
rect -1090 -1800 -1044 -1696
rect -966 -1708 -940 -1696
rect -744 -1596 -638 -1586
rect -744 -1638 -720 -1596
rect -662 -1638 -638 -1596
rect -966 -1800 -932 -1708
rect -1090 -1816 -932 -1800
rect -1072 -1994 -932 -1816
rect -744 -1858 -638 -1638
rect -744 -1900 -724 -1858
rect -666 -1900 -638 -1858
rect 1830 -1588 1914 -1568
rect 1830 -1630 1838 -1588
rect 1896 -1630 1914 -1588
rect 1830 -1806 1914 -1630
rect 2128 -1652 2256 -1498
rect 2128 -1734 2156 -1652
rect 1830 -1848 1836 -1806
rect 1894 -1848 1914 -1806
rect 1830 -1862 1914 -1848
rect 2120 -1758 2156 -1734
rect 2236 -1734 2256 -1652
rect 2236 -1758 2272 -1734
rect -744 -1908 -638 -1900
rect 1418 -1920 1550 -1918
rect 1322 -1940 1962 -1920
rect -1072 -2426 -1030 -1994
rect -960 -2426 -932 -1994
rect -1072 -2532 -932 -2426
rect -750 -1994 -108 -1974
rect -750 -2426 -712 -1994
rect -642 -2426 -108 -1994
rect -750 -2446 -108 -2426
rect -248 -2604 -108 -2446
rect 1322 -2372 1834 -1940
rect 1904 -2372 1962 -1940
rect 1322 -2392 1962 -2372
rect 2120 -1940 2272 -1758
rect 2120 -2372 2152 -1940
rect 2222 -2372 2272 -1940
rect 1322 -2562 1462 -2392
rect 2120 -2398 2272 -2372
rect -248 -2638 -232 -2604
rect -126 -2638 -108 -2604
rect -248 -2646 -108 -2638
rect -78 -2606 1288 -2586
rect 1322 -2596 1336 -2562
rect 1442 -2596 1462 -2562
rect 1322 -2606 1462 -2596
rect -78 -2608 1248 -2606
rect -78 -2648 164 -2608
rect -78 -2682 -72 -2648
rect -38 -2680 164 -2648
rect 234 -2640 1248 -2608
rect 1282 -2640 1288 -2606
rect 234 -2680 1288 -2640
rect -38 -2682 1288 -2680
rect -248 -2692 -110 -2684
rect -248 -2726 -232 -2692
rect -126 -2726 -110 -2692
rect -78 -2704 1288 -2682
rect 1324 -2650 1456 -2640
rect 1324 -2684 1336 -2650
rect 1442 -2684 1456 -2650
rect -248 -2752 -110 -2726
rect 1324 -2752 1456 -2684
rect 3106 -2651 3568 -2515
rect -584 -2764 1750 -2752
rect -584 -2770 1246 -2764
rect -584 -2796 -548 -2770
rect -512 -2796 1246 -2770
rect -584 -2856 -552 -2796
rect -494 -2800 1246 -2796
rect 1304 -2800 1370 -2764
rect 1428 -2800 1474 -2764
rect 1532 -2788 1750 -2764
rect 1532 -2800 1702 -2788
rect -494 -2804 1702 -2800
rect -494 -2840 -322 -2804
rect -264 -2806 -94 -2804
rect -264 -2840 -206 -2806
rect -494 -2842 -206 -2840
rect -148 -2840 -94 -2806
rect -36 -2824 1702 -2804
rect 1738 -2824 1750 -2788
rect -36 -2840 1750 -2824
rect -148 -2842 1750 -2840
rect -494 -2856 1750 -2842
rect -584 -2860 1750 -2856
rect -584 -2896 -546 -2860
rect -510 -2862 1750 -2860
rect -510 -2896 1702 -2862
rect -584 -2898 1702 -2896
rect 1738 -2898 1750 -2862
rect -584 -2918 1750 -2898
rect 3106 -2823 3245 -2651
rect 3438 -2823 3568 -2651
rect 272 -4327 734 -2918
rect 3106 -2960 3568 -2823
rect 272 -4499 411 -4327
rect 604 -4499 734 -4327
rect -1076 -4626 -614 -4604
rect -1076 -5058 -1030 -4626
rect -960 -5058 -712 -4626
rect -642 -5058 -614 -4626
rect 272 -4636 734 -4499
rect 1802 -4572 2264 -4550
rect 1802 -5004 1834 -4572
rect 1904 -5004 2152 -4572
rect 2222 -5004 2264 -4572
rect 1802 -5022 2264 -5004
rect -1076 -5076 -614 -5058
<< via1 >>
rect 411 534 604 706
rect -1294 272 -1240 324
rect -624 30 -572 84
rect -1044 -1800 -966 -1696
rect 2156 -1758 2236 -1652
rect 164 -2680 234 -2608
rect -552 -2806 -548 -2796
rect -548 -2806 -512 -2796
rect -512 -2806 -494 -2796
rect -552 -2856 -494 -2806
rect 3245 -2823 3438 -2651
rect 411 -4499 604 -4327
<< metal2 >>
rect 272 737 734 842
rect 272 504 380 737
rect 632 504 734 737
rect 272 397 734 504
rect -1316 324 -1234 330
rect -1316 320 -1294 324
rect -1318 260 -1306 320
rect -1240 272 -1234 324
rect -1246 260 -1234 272
rect -1318 252 -1234 260
rect -1316 248 -1234 252
rect -1374 84 -568 106
rect -1374 30 -624 84
rect -572 30 -568 84
rect -1374 0 -568 30
rect -1368 -120 -1246 0
rect -1364 -2760 -1248 -120
rect 2118 -1652 2284 -1636
rect -1096 -1680 -918 -1678
rect -1096 -1692 -916 -1680
rect -1096 -1696 -1034 -1692
rect -1096 -1800 -1044 -1696
rect -962 -1794 -916 -1692
rect 2118 -1758 2156 -1652
rect 2236 -1758 2284 -1652
rect 2118 -1792 2284 -1758
rect -966 -1800 -916 -1794
rect -1096 -1804 -916 -1800
rect -1096 -1810 -918 -1804
rect 3106 -2586 3568 -2515
rect 134 -2608 3568 -2586
rect 134 -2680 164 -2608
rect 234 -2620 3568 -2608
rect 234 -2680 3214 -2620
rect 134 -2706 3214 -2680
rect -1364 -2796 -474 -2760
rect -1364 -2856 -552 -2796
rect -494 -2856 -474 -2796
rect -1364 -2898 -474 -2856
rect 3106 -2853 3214 -2706
rect 3466 -2853 3568 -2620
rect -1364 -2900 -1248 -2898
rect 3106 -2960 3568 -2853
rect 272 -4296 734 -4191
rect 272 -4529 380 -4296
rect 632 -4529 734 -4296
rect 272 -4636 734 -4529
<< via2 >>
rect 380 706 632 737
rect 380 534 411 706
rect 411 534 604 706
rect 604 534 632 706
rect 380 504 632 534
rect -1306 272 -1294 320
rect -1294 272 -1246 320
rect -1306 260 -1246 272
rect -1034 -1696 -962 -1692
rect -1034 -1794 -966 -1696
rect -966 -1794 -962 -1696
rect 2156 -1758 2236 -1652
rect 164 -2680 234 -2608
rect 3214 -2651 3466 -2620
rect 3214 -2823 3245 -2651
rect 3245 -2823 3438 -2651
rect 3438 -2823 3466 -2651
rect 3214 -2853 3466 -2823
rect 380 -4327 632 -4296
rect 380 -4499 411 -4327
rect 411 -4499 604 -4327
rect 604 -4499 632 -4327
rect 380 -4529 632 -4499
<< metal3 >>
rect 272 760 734 842
rect 272 477 357 760
rect 656 477 734 760
rect 272 397 734 477
rect -1316 320 -1240 326
rect -1316 298 -1306 320
rect -1318 260 -1306 298
rect -1246 260 -1240 320
rect -1318 224 -1240 260
rect -1318 -2586 -1246 224
rect 2132 -1652 2264 -1636
rect -1088 -1692 -914 -1678
rect -1088 -1698 -1034 -1692
rect -1088 -1796 -1040 -1698
rect -962 -1794 -914 -1692
rect -964 -1796 -914 -1794
rect -1088 -1810 -914 -1796
rect 2132 -1758 2152 -1652
rect 2236 -1758 2264 -1652
rect 2132 -1800 2264 -1758
rect -1322 -2608 256 -2586
rect -1322 -2680 164 -2608
rect 234 -2680 256 -2608
rect -1322 -2706 256 -2680
rect 3106 -2597 3568 -2515
rect 3106 -2880 3191 -2597
rect 3490 -2880 3568 -2597
rect 3106 -2960 3568 -2880
rect 272 -4273 734 -4191
rect 272 -4556 357 -4273
rect 656 -4556 734 -4273
rect 272 -4636 734 -4556
<< via3 >>
rect 357 737 656 760
rect 357 504 380 737
rect 380 504 632 737
rect 632 504 656 737
rect 357 477 656 504
rect -1040 -1794 -1034 -1698
rect -1034 -1794 -964 -1698
rect -1040 -1796 -964 -1794
rect 2152 -1758 2156 -1652
rect 2156 -1758 2234 -1652
rect 3191 -2620 3490 -2597
rect 3191 -2853 3214 -2620
rect 3214 -2853 3466 -2620
rect 3466 -2853 3490 -2620
rect 3191 -2880 3490 -2853
rect 357 -4296 656 -4273
rect 357 -4529 380 -4296
rect 380 -4529 632 -4296
rect 632 -4529 656 -4296
rect 357 -4556 656 -4529
<< metal4 >>
rect 272 781 734 842
rect 272 452 333 781
rect 679 452 734 781
rect 272 397 734 452
rect 3106 -643 3568 -582
rect 3106 -804 3167 -643
rect -1077 -962 3167 -804
rect -3702 -1237 -3240 -1176
rect -3702 -1566 -3641 -1237
rect -3295 -1384 -3240 -1237
rect -3295 -1566 -2870 -1384
rect -3702 -1594 -2870 -1566
rect -3702 -1621 -3240 -1594
rect -1077 -1676 -914 -962
rect 3106 -972 3167 -962
rect 3513 -972 3568 -643
rect 3106 -1027 3568 -972
rect 3106 -1638 3568 -1610
rect -1620 -1698 -914 -1676
rect -1620 -1796 -1040 -1698
rect -964 -1796 -914 -1698
rect -1620 -1810 -914 -1796
rect 742 -1652 3568 -1638
rect 742 -1758 2152 -1652
rect 2234 -1665 3568 -1652
rect 2234 -1758 3167 -1665
rect 742 -1796 3167 -1758
rect 742 -2224 880 -1796
rect 3106 -1994 3167 -1796
rect 3513 -1994 3568 -1665
rect 3106 -2055 3568 -1994
rect -1506 -2358 886 -2224
rect 3106 -2576 3568 -2515
rect -3702 -2761 -3240 -2700
rect -3702 -3090 -3641 -2761
rect -3295 -2808 -3240 -2761
rect -3295 -3018 -2664 -2808
rect 3106 -2905 3167 -2576
rect 3513 -2905 3568 -2576
rect 3106 -2960 3568 -2905
rect -3295 -3090 -3240 -3018
rect -3702 -3145 -3240 -3090
rect 272 -4252 734 -4191
rect 272 -4581 333 -4252
rect 679 -4581 734 -4252
rect 272 -4636 734 -4581
<< via4 >>
rect 333 760 679 781
rect 333 477 357 760
rect 357 477 656 760
rect 656 477 679 760
rect 333 452 679 477
rect -3641 -1566 -3295 -1237
rect 3167 -972 3513 -643
rect 3167 -1994 3513 -1665
rect -3641 -3090 -3295 -2761
rect 3167 -2597 3513 -2576
rect 3167 -2880 3191 -2597
rect 3191 -2880 3490 -2597
rect 3490 -2880 3513 -2597
rect 3167 -2905 3513 -2880
rect 333 -4273 679 -4252
rect 333 -4556 357 -4273
rect 357 -4556 656 -4273
rect 656 -4556 679 -4273
rect 333 -4581 679 -4556
<< metal5 >>
rect 272 781 734 842
rect 272 452 333 781
rect 679 452 734 781
rect 272 397 734 452
rect 3106 -643 3568 -582
rect 3106 -972 3167 -643
rect 3513 -972 3568 -643
rect 3106 -1027 3568 -972
rect -3702 -1237 -3240 -1176
rect -3702 -1566 -3641 -1237
rect -3295 -1566 -3240 -1237
rect -3702 -1621 -3240 -1566
rect 3106 -1665 3568 -1610
rect 3106 -1994 3167 -1665
rect 3513 -1994 3568 -1665
rect 3106 -2055 3568 -1994
rect 3106 -2576 3568 -2515
rect -3702 -2761 -3240 -2700
rect -3702 -3090 -3641 -2761
rect -3295 -3090 -3240 -2761
rect 3106 -2905 3167 -2576
rect 3513 -2905 3568 -2576
rect 3106 -2960 3568 -2905
rect -3702 -3145 -3240 -3090
rect 272 -4252 734 -4191
rect 272 -4581 333 -4252
rect 679 -4581 734 -4252
rect 272 -4636 734 -4581
use sky130_fd_pr__cap_mim_m3_1_MCFBFU  sky130_fd_pr__cap_mim_m3_1_MCFBFU_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606253345
transform 1 0 -2212 0 1 -2784
box -786 -700 786 700
use sky130_fd_pr__cap_mim_m3_1_MCFBFU  sky130_fd_pr__cap_mim_m3_1_MCFBFU_1
timestamp 1606253345
transform 1 0 -2330 0 1 -1232
box -786 -700 786 700
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/CustomFlow/magic/Work-main/layouts/RingOscillator
timestamp 1606359646
transform 1 0 -634 0 1 56
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606097532
transform 0 1 252 -1 0 182
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_N92D86  sky130_fd_pr__nfet_01v8_N92D86_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606102148
transform 0 1 -179 -1 0 -2665
box -211 -275 211 275
use sky130_fd_pr__res_xhigh_po_0p35_RF56VW  sky130_fd_pr__res_xhigh_po_0p35_RF56VW_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606102148
transform 1 0 -836 0 1 -3526
box -360 -1698 360 1698
use sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ  sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606097532
transform 1 0 -371 0 1 -870
box -837 -798 837 798
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_1
timestamp 1606097532
transform 0 1 889 -1 0 183
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_N92D86  sky130_fd_pr__nfet_01v8_N92D86_1
timestamp 1606102148
transform 0 1 1389 -1 0 -2623
box -211 -275 211 275
use sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ  sky130_fd_pr__res_xhigh_po_0p35_YEQXSQ_1
timestamp 1606097532
transform 1 0 1555 0 1 -866
box -837 -798 837 798
use sky130_fd_pr__res_xhigh_po_0p35_RF56VW  sky130_fd_pr__res_xhigh_po_0p35_RF56VW_1
timestamp 1606102148
transform 1 0 2028 0 1 -3472
box -360 -1698 360 1698
<< labels >>
rlabel metal1 71 165 105 199 1 inv_out
rlabel metal1 556 342 590 376 1 Vdd
port 1 n
rlabel metal1 -1042 -1798 -962 -1690 1 VP
port 2 n
rlabel metal1 2154 -1760 2234 -1652 1 VN
port 3 n
rlabel metal1 532 -2660 590 -2606 1 C1
port 4 n
rlabel metal1 540 -2860 598 -2806 1 Gnd
port 5 n
rlabel via4 -3414 -1566 -3306 -1426 1 INP
port 6 n
rlabel metal4 -3180 -2974 -3072 -2834 1 INN
port 7 n
<< end >>
