magic
tech sky130A
magscale 1 2
timestamp 1606790247
<< nwell >>
rect -2760 4240 11100 4600
<< pwell >>
rect -2180 -3500 -2100 -3280
<< psubdiff >>
rect -2720 -3700 10560 -3680
rect -2720 -3740 -1620 -3700
rect 2800 -3740 10560 -3700
rect -2720 -3780 -2660 -3740
rect 10520 -3780 10560 -3740
rect -2720 -3820 -1620 -3780
rect 2800 -3820 10560 -3780
rect -2720 -3840 10560 -3820
<< nsubdiff >>
rect -2620 4460 10980 4480
rect -2620 4380 -2580 4460
rect 10920 4380 10980 4460
rect -2620 4360 10980 4380
<< psubdiffcont >>
rect -1620 -3740 2800 -3700
rect -2660 -3780 10520 -3740
rect -1620 -3820 2800 -3780
<< nsubdiffcont >>
rect -2580 4380 10920 4460
<< locali >>
rect -2620 4460 10980 4480
rect -2620 4380 -2580 4460
rect 10920 4380 10980 4460
rect 600 4360 10980 4380
rect -2720 -3700 10560 -3680
rect -2720 -3740 -1620 -3700
rect 2800 -3740 10560 -3700
rect -2720 -3780 -2660 -3740
rect 10520 -3780 10560 -3740
rect -2720 -3820 -1620 -3780
rect 2800 -3820 10560 -3780
rect -2720 -3840 10560 -3820
<< rlocali >>
rect -1760 -2200 -1740 -2080
<< viali >>
rect -2580 4380 10920 4460
rect -2380 4100 -2280 4140
rect -1900 4100 -1800 4140
rect -1460 4100 -1360 4140
rect -1000 4100 -900 4140
rect -540 4100 -440 4140
rect -80 4100 20 4140
rect 380 4100 480 4140
rect 2900 4100 3000 4140
rect 3360 4100 3460 4140
rect 3820 4100 3920 4140
rect 4280 4100 4380 4140
rect 4720 4100 4820 4140
rect 5200 4100 5300 4140
rect 5680 4100 5780 4140
rect 7920 4100 8020 4140
rect 8360 4100 8460 4140
rect 8820 4100 8920 4140
rect 9280 4100 9380 4140
rect 9740 4100 9840 4140
rect 10200 4100 10300 4140
rect 10660 4100 10760 4140
rect -2580 3620 -2540 3780
rect -1660 3620 -1620 3780
rect -740 3600 -700 3760
rect 160 3620 200 3780
rect 740 3620 780 3760
rect 2700 3600 2740 3760
rect 3620 3580 3660 3760
rect 4540 3580 4580 3760
rect 5460 3580 5500 3760
rect 6020 3620 6060 3760
rect 7600 3600 7640 3740
rect 7720 3600 7760 3720
rect 8640 3600 8680 3720
rect 9560 3600 9600 3720
rect 10480 3600 10520 3720
rect -2100 2960 -2060 3060
rect -1200 2960 -1160 3060
rect -280 2960 -240 3060
rect 640 2960 680 3060
rect 3160 2880 3200 3040
rect 4080 2880 4120 3040
rect 5000 2880 5040 3040
rect 5900 2880 5940 3040
rect 8160 2800 8200 2900
rect 9080 2800 9120 2900
rect 10000 2800 10040 2900
rect 10900 2800 10940 2900
rect 360 2580 460 2620
rect -1300 2300 -1220 2340
rect 4020 2300 4140 2340
rect 6900 2240 6960 2320
rect 1280 2100 1400 2140
rect 4040 2100 4160 2140
rect 6880 2100 7000 2140
rect 1280 2000 1400 2040
rect 4040 2000 4140 2040
rect 6880 2000 7020 2040
rect 2280 1820 2320 1920
rect 3360 1820 3400 1920
rect 4880 1820 4920 1920
rect 6160 1820 6200 1920
rect 2060 1720 2140 1760
rect 3540 1720 3700 1760
rect 6880 1720 7020 1760
rect 3520 1300 3680 1340
rect 4920 1280 5080 1320
rect 2060 900 2140 1180
rect 6880 1160 7020 1200
rect 6140 1020 6180 1060
rect 6580 900 6740 940
rect 7500 900 7660 940
rect -1340 680 -1300 860
rect 540 680 600 860
rect 1060 720 1100 840
rect 4940 820 5100 860
rect 6620 780 6700 820
rect 3280 660 3320 740
rect 5380 660 5420 740
rect 3700 540 3740 580
rect -1900 260 -1860 400
rect -1800 260 -1760 400
rect -20 240 20 380
rect 80 240 120 400
rect 2060 120 2140 500
rect 3660 440 3760 480
rect 5740 180 5820 220
rect -1620 40 -1460 100
rect 280 20 420 80
rect 2780 -720 2820 -580
rect 3700 -720 3740 -580
rect 4620 -700 4660 -560
rect 5540 -700 5580 -560
rect 6640 -720 6680 -560
rect 7560 -720 7600 -560
rect 8480 -700 8520 -540
rect 9400 -700 9440 -540
rect 3240 -1160 3280 -1060
rect 4160 -1160 4200 -1060
rect 5080 -1160 5120 -1060
rect 6000 -1160 6040 -1060
rect 6100 -1160 6140 -1080
rect 7100 -1160 7140 -1060
rect 8020 -1160 8060 -1060
rect 8940 -1160 8980 -1060
rect 9860 -1160 9900 -1060
rect 9960 -1140 10000 -1060
rect 2980 -1340 3100 -1300
rect 3460 -1340 3580 -1300
rect 3900 -1340 4020 -1300
rect 4360 -1340 4480 -1300
rect 4840 -1340 4960 -1300
rect 5280 -1340 5400 -1300
rect 5740 -1340 5860 -1300
rect 6840 -1340 6960 -1300
rect 7320 -1340 7440 -1300
rect 7760 -1340 7880 -1300
rect 8220 -1340 8340 -1300
rect 8680 -1340 8800 -1300
rect 9160 -1340 9280 -1300
rect 9620 -1340 9740 -1300
rect -1780 -2320 -1740 -2240
rect -860 -2320 -820 -2240
rect 60 -2320 100 -2240
rect 980 -2320 1020 -2240
rect 1900 -2320 1940 -2240
rect 2800 -2320 2840 -2240
rect 4960 -2360 5000 -2260
rect 5880 -2360 5920 -2260
rect 6800 -2360 6840 -2260
rect 7720 -2360 7760 -2260
rect 8640 -2360 8680 -2260
rect 9540 -2380 9580 -2280
rect 10460 -2380 10500 -2280
rect -2180 -3200 -2140 -3120
rect -2060 -3220 -2020 -3100
rect -1880 -3220 -1840 -3120
rect -1320 -3200 -1280 -3120
rect -400 -3200 -360 -3120
rect 520 -3200 560 -3120
rect 1440 -3200 1480 -3120
rect 2340 -3200 2380 -3120
rect 4860 -3200 4900 -3120
rect 5420 -3200 5460 -3120
rect 6340 -3200 6380 -3120
rect 7260 -3200 7300 -3120
rect 8160 -3200 8200 -3120
rect 9080 -3200 9120 -3120
rect 10000 -3200 10040 -3120
rect -2640 -3400 -2600 -3300
rect -2480 -3480 -2340 -3440
rect -1600 -3480 -1460 -3440
rect -1140 -3480 -1000 -3440
rect -680 -3480 -540 -3440
rect -260 -3480 -120 -3440
rect 220 -3480 360 -3440
rect 680 -3480 820 -3440
rect 1140 -3480 1280 -3440
rect 1600 -3480 1740 -3440
rect 2060 -3480 2200 -3440
rect 2540 -3480 2680 -3440
rect 5160 -3480 5280 -3440
rect 5620 -3480 5740 -3440
rect 6080 -3480 6200 -3440
rect 6540 -3480 6660 -3440
rect 7000 -3480 7120 -3440
rect 7440 -3480 7560 -3440
rect 7900 -3480 8020 -3440
rect 8360 -3480 8480 -3440
rect 8840 -3480 8960 -3440
rect 9280 -3480 9400 -3440
rect 9740 -3480 9860 -3440
rect 10200 -3480 10320 -3440
rect -2660 -3780 10520 -3740
<< metal1 >>
rect -2700 4460 11060 4520
rect -3480 4340 -3040 4420
rect -2700 4380 -2580 4460
rect 10920 4380 11060 4460
rect -2700 4340 11060 4380
rect -3480 4220 -3340 4340
rect -3160 4240 -2520 4340
rect -3160 4220 -3040 4240
rect -3480 4120 -3040 4220
rect -2620 3800 -2520 4240
rect -2420 4140 10920 4160
rect -2420 4100 -2380 4140
rect -2280 4100 -1900 4140
rect -1800 4100 -1460 4140
rect -1360 4100 -1000 4140
rect -900 4100 -540 4140
rect -440 4100 -80 4140
rect 20 4100 380 4140
rect 480 4100 2900 4140
rect 3000 4100 3360 4140
rect 3460 4100 3820 4140
rect 3920 4100 4280 4140
rect 4380 4100 4720 4140
rect 4820 4100 5200 4140
rect 5300 4100 5680 4140
rect 5780 4100 7920 4140
rect 8020 4100 8360 4140
rect 8460 4100 8820 4140
rect 8920 4100 9280 4140
rect 9380 4100 9740 4140
rect 9840 4100 10200 4140
rect 10300 4100 10660 4140
rect 10760 4100 10920 4140
rect -2420 4080 10920 4100
rect 2680 3800 5960 3820
rect -2620 3780 10560 3800
rect -2620 3620 -2580 3780
rect -2540 3620 -1660 3780
rect -1620 3760 160 3780
rect -1620 3620 -740 3760
rect -2620 3600 -740 3620
rect -700 3620 160 3760
rect 200 3760 10560 3780
rect 200 3620 740 3760
rect 780 3620 2700 3760
rect -700 3600 2700 3620
rect 2740 3600 3620 3760
rect -2620 3580 3620 3600
rect 3660 3580 4540 3760
rect 4580 3580 5460 3760
rect 5500 3620 6020 3760
rect 6060 3740 10560 3760
rect 6060 3620 7600 3740
rect 5500 3600 7600 3620
rect 7640 3720 10560 3740
rect 7640 3600 7720 3720
rect 7760 3600 8640 3720
rect 8680 3600 9560 3720
rect 9600 3600 10480 3720
rect 10520 3600 10560 3720
rect 5500 3580 10560 3600
rect -2620 3540 10560 3580
rect -2120 3120 700 3140
rect -2120 3060 1480 3120
rect -2120 2960 -2100 3060
rect -2060 2960 -1200 3060
rect -1160 2960 -280 3060
rect -240 2960 640 3060
rect 680 2960 1480 3060
rect -2120 2880 1480 2960
rect 320 2620 480 2640
rect 320 2580 360 2620
rect 460 2580 480 2620
rect -1340 2360 -1160 2380
rect -1340 2280 -1320 2360
rect -1220 2280 -1160 2360
rect -1340 2220 -1160 2280
rect -1340 880 -1260 2220
rect 320 1760 480 2580
rect 1200 2140 1480 2880
rect 3140 3040 5960 3200
rect 3140 2880 3160 3040
rect 3200 2880 4080 3040
rect 4120 2880 5000 3040
rect 5040 2880 5900 3040
rect 5940 2880 5960 3040
rect 3140 2840 5960 2880
rect 6800 2900 10960 3000
rect 1200 2100 1280 2140
rect 1400 2100 1480 2140
rect 1200 2040 1480 2100
rect 1200 2000 1280 2040
rect 1400 2000 1480 2040
rect 1200 1980 1480 2000
rect 3980 2360 4200 2840
rect 4180 2260 4200 2360
rect 3980 2140 4200 2260
rect 3980 2100 4040 2140
rect 4160 2100 4200 2140
rect 3980 2040 4200 2100
rect 3980 2000 4040 2040
rect 4140 2000 4200 2040
rect 3980 1980 4200 2000
rect 6800 2800 8160 2900
rect 8200 2800 9080 2900
rect 9120 2800 10000 2900
rect 10040 2800 10900 2900
rect 10940 2800 10960 2900
rect 6800 2720 10960 2800
rect 6800 2360 7100 2720
rect 6800 2200 6820 2360
rect 7040 2200 7100 2360
rect 6800 2140 7100 2200
rect 6800 2100 6880 2140
rect 7000 2100 7100 2140
rect 6800 2040 7100 2100
rect 6800 2000 6880 2040
rect 7020 2000 7100 2040
rect 6800 1980 7100 2000
rect 2260 1920 3420 1980
rect 2260 1820 2280 1920
rect 2320 1820 3360 1920
rect 3400 1820 3420 1920
rect 2260 1780 3420 1820
rect 4860 1920 6220 1980
rect 4860 1820 4880 1920
rect 4920 1820 6160 1920
rect 6200 1820 6220 1920
rect 4860 1780 6220 1820
rect 2020 1760 2180 1780
rect 320 1720 2060 1760
rect 2140 1720 2180 1760
rect 320 1680 2180 1720
rect 2020 1180 2180 1680
rect 2020 900 2060 1180
rect 2140 900 2180 1180
rect -1360 860 -1260 880
rect -1360 680 -1340 860
rect -1300 700 -1260 860
rect 500 860 1180 880
rect 2020 860 2180 900
rect -1300 680 -1280 700
rect -1360 660 -1280 680
rect 500 680 540 860
rect 600 700 980 860
rect 600 680 1180 700
rect 500 660 1180 680
rect 2020 500 2200 540
rect -1800 440 -1740 500
rect -1920 400 -1740 440
rect 60 420 120 500
rect -1920 260 -1900 400
rect -1860 260 -1800 400
rect -1760 260 -1740 400
rect -1920 240 -1740 260
rect -1800 -2200 -1740 240
rect -40 400 140 420
rect -40 380 80 400
rect -40 240 -20 380
rect 20 240 80 380
rect 120 240 140 400
rect -40 220 140 240
rect -1640 100 -1440 120
rect -1640 40 -1620 100
rect -1460 40 -1440 100
rect -1640 -120 -1440 40
rect -920 -80 -480 0
rect -920 -120 -780 -80
rect -1640 -200 -780 -120
rect -600 -200 -480 -80
rect -1640 -240 -480 -200
rect -1640 -320 -1440 -240
rect -920 -300 -480 -240
rect 60 -2200 120 220
rect 2020 120 2060 500
rect 2140 120 2200 500
rect 2020 100 2180 120
rect 240 80 440 100
rect 240 20 280 80
rect 420 20 440 80
rect 240 -120 440 20
rect 840 -120 1280 -40
rect 240 -240 980 -120
rect 1160 -240 1280 -120
rect 240 -320 440 -240
rect 840 -340 1280 -240
rect 2060 -1580 2140 100
rect 2300 -1580 2440 1780
rect 3460 1760 3780 1780
rect 4880 1760 6220 1780
rect 6800 1760 7080 1780
rect 3460 1720 3540 1760
rect 3700 1720 3780 1760
rect 3460 1340 3780 1720
rect 6800 1720 6880 1760
rect 7020 1720 7080 1760
rect 6800 1500 7080 1720
rect 8520 1500 8960 1580
rect 6800 1380 8660 1500
rect 8840 1380 8960 1500
rect 6800 1360 8960 1380
rect 3460 1300 3520 1340
rect 3680 1300 3780 1340
rect 3460 1260 3780 1300
rect 4860 1320 5840 1340
rect 4860 1280 4920 1320
rect 5080 1280 5840 1320
rect 4860 1260 5840 1280
rect 3500 1080 3700 1260
rect 3260 1020 3700 1080
rect 3260 740 3340 1020
rect 4860 860 5180 1260
rect 4860 820 4940 860
rect 5100 820 5180 860
rect 4860 800 5180 820
rect 3260 660 3280 740
rect 3320 660 3340 740
rect 3260 620 3340 660
rect 5360 740 5440 760
rect 5360 620 5440 660
rect 3680 580 3760 600
rect 3680 540 3700 580
rect 3740 540 3760 580
rect 3680 500 3760 540
rect 3620 480 3800 500
rect 3620 440 3660 480
rect 3760 440 3800 480
rect 3620 420 3800 440
rect 3700 -500 3740 420
rect 5720 220 5840 1260
rect 6800 1200 7080 1360
rect 8520 1280 8960 1360
rect 6800 1160 6880 1200
rect 7020 1160 7080 1200
rect 6800 1140 7080 1160
rect 6100 1000 6120 1080
rect 6200 1000 6220 1080
rect 6560 940 6760 960
rect 6560 900 6580 940
rect 6740 900 6760 940
rect 6560 880 6760 900
rect 7460 940 7680 960
rect 7460 900 7500 940
rect 7660 900 7680 940
rect 7460 880 7680 900
rect 6640 840 6680 880
rect 6600 820 6720 840
rect 6600 780 6620 820
rect 6700 780 6720 820
rect 6600 760 6720 780
rect 5720 180 5740 220
rect 5820 180 5840 220
rect 5720 160 5840 180
rect 6640 -500 6680 760
rect 7560 -500 7600 880
rect 2760 -560 5600 -500
rect 2760 -580 4620 -560
rect 2760 -720 2780 -580
rect 2820 -720 3700 -580
rect 3740 -700 4620 -580
rect 4660 -700 5540 -560
rect 5580 -700 5600 -560
rect 3740 -720 5600 -700
rect 2760 -760 5600 -720
rect 6620 -540 9460 -500
rect 6620 -560 8480 -540
rect 6620 -720 6640 -560
rect 6680 -720 7560 -560
rect 7600 -700 8480 -560
rect 8520 -700 9400 -540
rect 9440 -700 9460 -540
rect 7600 -720 9460 -700
rect 6620 -760 9460 -720
rect 6620 -780 6700 -760
rect 3220 -1060 10920 -1020
rect 3220 -1160 3240 -1060
rect 3280 -1160 4160 -1060
rect 4200 -1160 5080 -1060
rect 5120 -1160 6000 -1060
rect 6040 -1080 7100 -1060
rect 6040 -1160 6100 -1080
rect 6140 -1160 7100 -1080
rect 7140 -1160 8020 -1060
rect 8060 -1160 8940 -1060
rect 8980 -1160 9860 -1060
rect 9900 -1140 9960 -1060
rect 10000 -1140 10920 -1060
rect 9900 -1160 10920 -1140
rect 3220 -1180 10920 -1160
rect 2840 -1300 9840 -1260
rect 2840 -1340 2980 -1300
rect 3100 -1340 3460 -1300
rect 3580 -1340 3900 -1300
rect 4020 -1340 4360 -1300
rect 4480 -1340 4840 -1300
rect 4960 -1340 5280 -1300
rect 5400 -1340 5740 -1300
rect 5860 -1340 6840 -1300
rect 6960 -1340 7320 -1300
rect 7440 -1340 7760 -1300
rect 7880 -1340 8220 -1300
rect 8340 -1340 8680 -1300
rect 8800 -1340 9160 -1300
rect 9280 -1340 9620 -1300
rect 9740 -1340 9840 -1300
rect 2840 -1360 9840 -1340
rect 2060 -1740 4000 -1580
rect 3820 -2180 4000 -1740
rect -1800 -2240 2860 -2200
rect -1800 -2320 -1780 -2240
rect -1740 -2320 -860 -2240
rect -820 -2320 60 -2240
rect 100 -2320 980 -2240
rect 1020 -2320 1900 -2240
rect 1940 -2320 2800 -2240
rect 2840 -2320 2860 -2240
rect -1800 -2380 2860 -2320
rect 3820 -2260 10520 -2180
rect 3820 -2360 4960 -2260
rect 5000 -2360 5880 -2260
rect 5920 -2360 6800 -2260
rect 6840 -2360 7720 -2260
rect 7760 -2360 8640 -2260
rect 8680 -2280 10520 -2260
rect 8680 -2360 9540 -2280
rect 3820 -2380 9540 -2360
rect 9580 -2380 10460 -2280
rect 10500 -2380 10520 -2280
rect 3820 -2440 10520 -2380
rect -2080 -3100 -2000 -3080
rect -1920 -3100 -1840 -3080
rect 10720 -3100 10920 -1180
rect -2200 -3120 -2060 -3100
rect -3520 -3260 -3080 -3180
rect -2200 -3200 -2180 -3120
rect -2140 -3200 -2060 -3120
rect -2200 -3220 -2060 -3200
rect -2020 -3120 10920 -3100
rect -2020 -3220 -1880 -3120
rect -1840 -3200 -1320 -3120
rect -1280 -3200 -400 -3120
rect -360 -3200 520 -3120
rect 560 -3200 1440 -3120
rect 1480 -3200 2340 -3120
rect 2380 -3200 4860 -3120
rect 4900 -3200 5420 -3120
rect 5460 -3200 6340 -3120
rect 6380 -3200 7260 -3120
rect 7300 -3200 8160 -3120
rect 8200 -3200 9080 -3120
rect 9120 -3200 10000 -3120
rect 10040 -3200 10920 -3120
rect -1840 -3220 10920 -3200
rect -2080 -3240 -2000 -3220
rect -1920 -3240 -1820 -3220
rect -3520 -3380 -3380 -3260
rect -3200 -3280 -3080 -3260
rect -3200 -3300 -2580 -3280
rect -3200 -3380 -2640 -3300
rect -3520 -3400 -2640 -3380
rect -2600 -3400 -2580 -3300
rect -3520 -3420 -2580 -3400
rect -1320 -3420 -1280 -3220
rect -400 -3420 -360 -3220
rect -3520 -3480 -3080 -3420
rect -2660 -3440 10460 -3420
rect -2660 -3480 -2480 -3440
rect -2340 -3480 -1600 -3440
rect -1460 -3480 -1140 -3440
rect -1000 -3480 -680 -3440
rect -540 -3480 -260 -3440
rect -120 -3480 220 -3440
rect 360 -3480 680 -3440
rect 820 -3480 1140 -3440
rect 1280 -3480 1600 -3440
rect 1740 -3480 2060 -3440
rect 2200 -3480 2540 -3440
rect 2680 -3480 5160 -3440
rect 5280 -3480 5620 -3440
rect 5740 -3480 6080 -3440
rect 6200 -3480 6540 -3440
rect 6660 -3480 7000 -3440
rect 7120 -3480 7440 -3440
rect 7560 -3480 7900 -3440
rect 8020 -3480 8360 -3440
rect 8480 -3480 8840 -3440
rect 8960 -3480 9280 -3440
rect 9400 -3480 9740 -3440
rect 9860 -3480 10200 -3440
rect 10320 -3480 10460 -3440
rect -2660 -3494 10460 -3480
rect -2660 -3498 -404 -3494
rect -2660 -3500 -1328 -3498
rect -1272 -3500 -404 -3498
rect -348 -3500 10460 -3494
rect -400 -3620 -360 -3618
rect -2780 -3622 -1328 -3620
rect -1272 -3622 10640 -3620
rect -2780 -3740 10640 -3622
rect -2780 -3780 -2660 -3740
rect 10520 -3780 10640 -3740
rect -2780 -3880 10640 -3780
rect -1820 -4060 -1700 -3880
rect -2000 -4140 -1560 -4060
rect -2000 -4260 -1860 -4140
rect -1680 -4260 -1560 -4140
rect -2000 -4360 -1560 -4260
<< via1 >>
rect -3340 4220 -3160 4340
rect -1320 2340 -1220 2360
rect -1320 2300 -1300 2340
rect -1300 2300 -1220 2340
rect -1320 2280 -1220 2300
rect 3980 2340 4180 2360
rect 3980 2300 4020 2340
rect 4020 2300 4140 2340
rect 4140 2300 4180 2340
rect 3980 2260 4180 2300
rect 6820 2320 7040 2360
rect 6820 2240 6900 2320
rect 6900 2240 6960 2320
rect 6960 2240 7040 2320
rect 6820 2200 7040 2240
rect 980 840 1180 860
rect 980 720 1060 840
rect 1060 720 1100 840
rect 1100 720 1180 840
rect 980 700 1180 720
rect -780 -200 -600 -80
rect 980 -240 1160 -120
rect 8660 1380 8840 1500
rect 5360 660 5380 740
rect 5380 660 5420 740
rect 5420 660 5440 740
rect 6120 1060 6200 1080
rect 6120 1020 6140 1060
rect 6140 1020 6180 1060
rect 6180 1020 6200 1060
rect 6120 1000 6200 1020
rect -3380 -3380 -3200 -3260
rect -1860 -4260 -1680 -4140
<< metal2 >>
rect -3500 4360 -3000 4460
rect -3500 4200 -3380 4360
rect -3120 4200 -3000 4360
rect -3500 4080 -3000 4200
rect -1340 2360 4200 2380
rect -1340 2280 -1320 2360
rect -1220 2280 3980 2360
rect -1340 2260 3980 2280
rect 4180 2260 4200 2360
rect -1340 2220 4200 2260
rect 5680 2360 7100 2380
rect 5680 2200 6820 2360
rect 7040 2200 7100 2360
rect 5680 1540 5900 2200
rect 980 1340 5900 1540
rect 8500 1520 9000 1620
rect 8500 1360 8620 1520
rect 8880 1360 9000 1520
rect 980 860 1180 1340
rect 8500 1240 9000 1360
rect 6100 1080 6220 1120
rect 6100 1000 6120 1080
rect 6200 1000 6220 1080
rect 6100 920 6220 1000
rect 6120 780 6200 920
rect 980 680 1180 700
rect 5340 740 6200 780
rect 5340 660 5360 740
rect 5440 660 6200 740
rect 5340 620 6200 660
rect -940 -60 -440 40
rect -940 -220 -820 -60
rect -560 -220 -440 -60
rect -940 -340 -440 -220
rect 820 -100 1320 0
rect 820 -260 940 -100
rect 1200 -260 1320 -100
rect 820 -380 1320 -260
rect -3540 -3240 -3040 -3140
rect -3540 -3400 -3420 -3240
rect -3160 -3400 -3040 -3240
rect -3540 -3520 -3040 -3400
rect -2020 -4120 -1520 -4020
rect -2020 -4280 -1900 -4120
rect -1640 -4280 -1520 -4120
rect -2020 -4400 -1520 -4280
<< via2 >>
rect -3380 4340 -3120 4360
rect -3380 4220 -3340 4340
rect -3340 4220 -3160 4340
rect -3160 4220 -3120 4340
rect -3380 4200 -3120 4220
rect 8620 1500 8880 1520
rect 8620 1380 8660 1500
rect 8660 1380 8840 1500
rect 8840 1380 8880 1500
rect 8620 1360 8880 1380
rect -820 -80 -560 -60
rect -820 -200 -780 -80
rect -780 -200 -600 -80
rect -600 -200 -560 -80
rect -820 -220 -560 -200
rect 940 -120 1200 -100
rect 940 -240 980 -120
rect 980 -240 1160 -120
rect 1160 -240 1200 -120
rect 940 -260 1200 -240
rect -3420 -3260 -3160 -3240
rect -3420 -3380 -3380 -3260
rect -3380 -3380 -3200 -3260
rect -3200 -3380 -3160 -3260
rect -3420 -3400 -3160 -3380
rect -1900 -4140 -1640 -4120
rect -1900 -4260 -1860 -4140
rect -1860 -4260 -1680 -4140
rect -1680 -4260 -1640 -4140
rect -1900 -4280 -1640 -4260
<< metal3 >>
rect -3520 4380 -2980 4460
rect -3520 4160 -3400 4380
rect -3100 4160 -2980 4380
rect -3520 4060 -2980 4160
rect 8480 1540 9020 1620
rect 8480 1320 8600 1540
rect 8900 1320 9020 1540
rect 8480 1220 9020 1320
rect -960 -40 -420 40
rect -960 -260 -840 -40
rect -540 -260 -420 -40
rect -960 -360 -420 -260
rect 800 -80 1340 0
rect 800 -300 920 -80
rect 1220 -300 1340 -80
rect 800 -400 1340 -300
rect -3560 -3220 -3020 -3140
rect -3560 -3440 -3440 -3220
rect -3140 -3440 -3020 -3220
rect -3560 -3540 -3020 -3440
rect -2040 -4100 -1500 -4020
rect -2040 -4320 -1920 -4100
rect -1620 -4320 -1500 -4100
rect -2040 -4420 -1500 -4320
<< via3 >>
rect -3400 4360 -3100 4380
rect -3400 4200 -3380 4360
rect -3380 4200 -3120 4360
rect -3120 4200 -3100 4360
rect -3400 4160 -3100 4200
rect 8600 1520 8900 1540
rect 8600 1360 8620 1520
rect 8620 1360 8880 1520
rect 8880 1360 8900 1520
rect 8600 1320 8900 1360
rect -840 -60 -540 -40
rect -840 -220 -820 -60
rect -820 -220 -560 -60
rect -560 -220 -540 -60
rect -840 -260 -540 -220
rect 920 -100 1220 -80
rect 920 -260 940 -100
rect 940 -260 1200 -100
rect 1200 -260 1220 -100
rect 920 -300 1220 -260
rect -3440 -3240 -3140 -3220
rect -3440 -3400 -3420 -3240
rect -3420 -3400 -3160 -3240
rect -3160 -3400 -3140 -3240
rect -3440 -3440 -3140 -3400
rect -1920 -4120 -1620 -4100
rect -1920 -4280 -1900 -4120
rect -1900 -4280 -1640 -4120
rect -1640 -4280 -1620 -4120
rect -1920 -4320 -1620 -4280
<< metal4 >>
rect -3540 4400 -2940 4480
rect -3540 4140 -3420 4400
rect -3080 4140 -2940 4400
rect -3540 4040 -2940 4140
rect 8460 1560 9060 1640
rect 8460 1300 8580 1560
rect 8920 1300 9060 1560
rect 8460 1200 9060 1300
rect -980 -20 -380 60
rect -980 -280 -860 -20
rect -520 -280 -380 -20
rect -980 -380 -380 -280
rect 780 -60 1380 20
rect 780 -320 900 -60
rect 1240 -320 1380 -60
rect 780 -420 1380 -320
rect -3580 -3200 -2980 -3120
rect -3580 -3460 -3460 -3200
rect -3120 -3460 -2980 -3200
rect -3580 -3560 -2980 -3460
rect -2060 -4080 -1460 -4000
rect -2060 -4340 -1940 -4080
rect -1600 -4340 -1460 -4080
rect -2060 -4440 -1460 -4340
<< via4 >>
rect -3420 4380 -3080 4400
rect -3420 4160 -3400 4380
rect -3400 4160 -3100 4380
rect -3100 4160 -3080 4380
rect -3420 4140 -3080 4160
rect 8580 1540 8920 1560
rect 8580 1320 8600 1540
rect 8600 1320 8900 1540
rect 8900 1320 8920 1540
rect 8580 1300 8920 1320
rect -860 -40 -520 -20
rect -860 -260 -840 -40
rect -840 -260 -540 -40
rect -540 -260 -520 -40
rect -860 -280 -520 -260
rect 900 -80 1240 -60
rect 900 -300 920 -80
rect 920 -300 1220 -80
rect 1220 -300 1240 -80
rect 900 -320 1240 -300
rect -3460 -3220 -3120 -3200
rect -3460 -3440 -3440 -3220
rect -3440 -3440 -3140 -3220
rect -3140 -3440 -3120 -3220
rect -3460 -3460 -3120 -3440
rect -1940 -4100 -1600 -4080
rect -1940 -4320 -1920 -4100
rect -1920 -4320 -1620 -4100
rect -1620 -4320 -1600 -4100
rect -1940 -4340 -1600 -4320
<< metal5 >>
rect -3560 4400 -2920 4500
rect -3560 4140 -3420 4400
rect -3080 4140 -2920 4400
rect -3560 4020 -2920 4140
rect 8440 1560 9080 1660
rect 8440 1300 8580 1560
rect 8920 1300 9080 1560
rect 8440 1180 9080 1300
rect -1000 -20 -360 80
rect -1000 -280 -860 -20
rect -520 -280 -360 -20
rect -1000 -400 -360 -280
rect 760 -60 1400 40
rect 760 -320 900 -60
rect 1240 -320 1400 -60
rect 760 -440 1400 -320
rect -3600 -3200 -2960 -3100
rect -3600 -3460 -3460 -3200
rect -3120 -3460 -2960 -3200
rect -3600 -3580 -2960 -3460
rect -2080 -4080 -1440 -3980
rect -2080 -4340 -1940 -4080
rect -1600 -4340 -1440 -4080
rect -2080 -4460 -1440 -4340
use sky130_fd_pr__nfet_01v8_lvt_4oweb9  sky130_fd_pr__nfet_01v8_lvt_4oweb9_0 arsalan
timestamp 1606578544
transform 1 0 -2384 0 1 -2710
box -396 -910 396 910
use sky130_fd_pr__nfet_01v8_lvt_goblxe  sky130_fd_pr__nfet_01v8_lvt_goblxe_0 arsalan
timestamp 1606471058
transform 1 0 537 0 1 -2710
box -2457 -910 2457 910
use sky130_fd_pr__nfet_01v8_lvt_6vyjkp  sky130_fd_pr__nfet_01v8_lvt_6vyjkp_0 arsalan
timestamp 1606471058
transform 1 0 7735 0 1 -2710
box -2915 -910 2915 910
use sky130_fd_pr__nfet_01v8_im9uye  sky130_fd_pr__nfet_01v8_im9uye_0 arsalan
timestamp 1606578544
transform 1 0 4410 0 1 -570
box -1770 -910 1770 910
use sky130_fd_pr__nfet_01v8_lvt_jzhy8l  sky130_fd_pr__nfet_01v8_lvt_jzhy8l_0 arsalan
timestamp 1606637863
transform 1 0 336 0 1 610
box -396 -710 396 710
use sky130_fd_pr__nfet_01v8_lvt_v5975p  sky130_fd_pr__nfet_01v8_lvt_v5975p_0 arsalan
timestamp 1606637863
transform 1 0 -1544 0 1 630
box -396 -710 396 710
use sky130_fd_pr__res_high_po_0p35_rfxuin  sky130_fd_pr__res_high_po_0p35_rfxuin_0 arsalan
timestamp 1606578544
transform 1 0 2101 0 1 689
box -201 -729 201 729
use sky130_fd_pr__nfet_01v8_cvwdxd  sky130_fd_pr__nfet_01v8_cvwdxd_0 arsalan
timestamp 1606578544
transform 1 0 8270 0 1 -570
box -1770 -910 1770 910
use sky130_fd_pr__pfet_01v8_lvt_2yzqpc  sky130_fd_pr__pfet_01v8_lvt_2yzqpc_0 arsalan
timestamp 1606471058
transform 0 1 1539 -1 0 1876
box -296 -919 296 919
use sky130_fd_pr__res_high_po_0p35_1pdy3p  sky130_fd_pr__res_high_po_0p35_1pdy3p_0 arsalan
timestamp 1606578544
transform 0 1 4337 -1 0 1301
box -201 -1057 201 1057
use sky130_fd_pr__nfet_01v8_lvt_u5ko20  sky130_fd_pr__nfet_01v8_lvt_u5ko20_0 arsalan
timestamp 1606578544
transform 0 1 4350 -1 0 696
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_lvt_m4eqfc  sky130_fd_pr__pfet_01v8_lvt_m4eqfc_0 arsalan
timestamp 1606578544
transform 0 1 6939 -1 0 1876
box -296 -919 296 919
use sky130_fd_pr__pfet_01v8_lvt_3xc4q5  sky130_fd_pr__pfet_01v8_lvt_3xc4q5_0 arsalan
timestamp 1606578544
transform 0 1 4139 -1 0 1876
box -296 -919 296 919
use sky130_fd_pr__nfet_01v8_lvt_gh6pom  sky130_fd_pr__nfet_01v8_lvt_gh6pom_0 arsalan
timestamp 1606578544
transform 0 1 7217 -1 0 1043
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_ekly11  sky130_fd_pr__pfet_01v8_ekly11_0 arsalan
timestamp 1606471058
transform 1 0 4330 0 1 3359
box -1770 -919 1770 919
use sky130_fd_pr__pfet_01v8_knu0r2  sky130_fd_pr__pfet_01v8_knu0r2_0 arsalan
timestamp 1606471058
transform 1 0 -950 0 1 3359
box -1770 -919 1770 919
use sky130_fd_pr__pfet_01v8_4yvul7  sky130_fd_pr__pfet_01v8_4yvul7_0 arsalan
timestamp 1606471058
transform 1 0 9330 0 1 3359
box -1770 -919 1770 919
<< labels >>
rlabel metal1 -2600 4260 -2540 4320 1 VDD
port 1 n
rlabel metal1 6860 1360 7060 1480 1 VOUT
port 2 n
rlabel metal1 -1580 -220 -1480 -120 1 VINP
port 3 n
rlabel metal1 300 -240 380 -120 1 VINN
port 4 n
rlabel metal1 -2880 -3380 -2800 -3320 1 IBP
port 5 n
rlabel metal1 -1800 -3840 -1700 -3680 1 VSS
port 6 n
<< end >>
