magic
tech sky130A
magscale 1 2
timestamp 1606621314
<< pwell >>
rect 1274 36 2630 1758
rect 272 -746 1150 12
rect 1274 -58 3248 36
rect 1570 -436 2096 -114
rect 1570 -437 1978 -436
rect 1570 -440 1930 -437
rect 1573 -442 1930 -440
rect 1573 -443 1978 -442
rect 1984 -443 2096 -436
rect 1573 -447 2096 -443
rect 1570 -644 2096 -447
rect 2370 -375 3248 -58
rect 2370 -709 2386 -375
rect 2370 -722 3248 -709
<< poly >>
rect 1386 -298 1482 -238
rect 1988 -298 2084 -238
rect 1372 -520 1537 -454
rect 1970 -514 2137 -448
<< locali >>
rect 186 2038 3244 2060
rect 186 1972 242 2038
rect 314 2036 2458 2038
rect 314 2032 2018 2036
rect 314 1972 552 2032
rect 186 1966 552 1972
rect 624 2026 1344 2032
rect 624 1966 868 2026
rect 186 1960 868 1966
rect 940 1966 1344 2026
rect 1416 1970 2018 2032
rect 2090 1972 2458 2036
rect 2530 1972 2752 2038
rect 2824 1972 3054 2038
rect 3126 1972 3244 2038
rect 2090 1970 3244 1972
rect 1416 1966 3244 1970
rect 940 1960 3244 1966
rect 186 1936 3244 1960
rect 1372 -476 1537 -470
rect 1372 -514 1377 -476
rect 1532 -514 1537 -476
rect 1970 -474 2137 -464
rect 1970 -510 1974 -474
rect 2132 -510 2137 -474
rect 1970 -514 2137 -510
rect 1372 -520 1537 -514
<< rlocali >>
rect 2238 -896 2242 -862
rect 2238 -898 2276 -896
<< viali >>
rect 242 1972 314 2038
rect 552 1966 624 2032
rect 868 1960 940 2026
rect 1344 1966 1416 2032
rect 2018 1970 2090 2036
rect 2458 1972 2530 2038
rect 2752 1972 2824 2038
rect 3054 1972 3126 2038
rect 113 1165 183 1597
rect 431 1165 501 1597
rect 749 1165 819 1597
rect 1067 1165 1137 1597
rect 2316 1160 2386 1592
rect 2634 1160 2704 1592
rect 2952 1160 3022 1592
rect 3270 1160 3340 1592
rect 113 113 183 545
rect 431 113 501 545
rect 749 113 819 545
rect 1067 113 1137 545
rect 2316 108 2386 540
rect 2634 108 2704 540
rect 2952 108 3022 540
rect 3270 108 3340 540
rect 240 -16 312 20
rect 608 -16 680 20
rect 920 -16 992 20
rect 2282 -22 3374 12
rect 1222 -408 1258 -346
rect 1338 -422 1372 -336
rect 1434 -422 1468 -336
rect 1530 -422 1564 -336
rect 1644 -408 1680 -346
rect 1826 -414 1862 -352
rect 1940 -420 1974 -334
rect 2036 -420 2070 -334
rect 2132 -420 2166 -334
rect 2246 -404 2282 -342
rect 1377 -514 1532 -476
rect 1974 -510 2132 -474
rect 490 -908 1466 -874
rect 2242 -896 2280 -860
rect 406 -1304 440 -936
rect 1516 -1304 1550 -936
rect 1968 -1292 2002 -924
rect 934 -1366 1070 -1332
rect 2494 -1354 2626 -1320
rect 400 -1480 1556 -1446
rect 1962 -1468 3118 -1434
<< metal1 >>
rect 94 2106 3230 2114
rect 94 2057 3360 2106
rect 94 1921 150 2057
rect 3286 1921 3360 2057
rect 94 1888 3360 1921
rect 94 1597 206 1888
rect 94 1165 113 1597
rect 183 1165 206 1597
rect 94 1142 206 1165
rect 404 1597 842 1626
rect 404 1165 431 1597
rect 501 1165 749 1597
rect 819 1165 842 1597
rect 404 1136 842 1165
rect 1044 1597 1474 1622
rect 1044 1165 1067 1597
rect 1137 1538 1474 1597
rect 1137 1197 1196 1538
rect 1392 1197 1474 1538
rect 1137 1165 1474 1197
rect 1044 1148 1474 1165
rect 88 545 524 564
rect 88 113 113 545
rect 183 113 431 545
rect 501 113 524 545
rect 88 90 524 113
rect 732 545 1154 560
rect 732 113 749 545
rect 819 113 1067 545
rect 1137 113 1154 545
rect 732 102 1154 113
rect 964 28 1206 30
rect 68 20 1206 28
rect 68 -16 240 20
rect 312 -16 608 20
rect 680 -16 920 20
rect 992 -16 1206 20
rect 68 -28 1206 -16
rect 224 -1402 350 -28
rect 1218 -318 1378 -316
rect 1212 -336 1378 -318
rect 1212 -346 1338 -336
rect 1212 -408 1222 -346
rect 1258 -408 1338 -346
rect 1212 -422 1338 -408
rect 1372 -422 1378 -336
rect 1212 -440 1378 -422
rect 1428 -336 1474 1148
rect 2004 1592 2414 1610
rect 2004 1546 2316 1592
rect 2004 1193 2056 1546
rect 2249 1193 2316 1546
rect 2004 1160 2316 1193
rect 2386 1160 2414 1592
rect 2004 1142 2414 1160
rect 2616 1592 3040 1616
rect 2616 1160 2634 1592
rect 2704 1160 2952 1592
rect 3022 1160 3040 1592
rect 2616 1142 3040 1160
rect 3254 1592 3360 1888
rect 3254 1160 3270 1592
rect 3340 1160 3360 1592
rect 3254 1144 3360 1160
rect 1822 -316 1982 -314
rect 1816 -320 1982 -316
rect 1428 -422 1434 -336
rect 1468 -422 1474 -336
rect 1428 -434 1474 -422
rect 1524 -334 1982 -320
rect 1524 -336 1940 -334
rect 1524 -422 1530 -336
rect 1564 -346 1940 -336
rect 1564 -408 1644 -346
rect 1680 -352 1940 -346
rect 1680 -408 1826 -352
rect 1564 -414 1826 -408
rect 1862 -414 1940 -352
rect 1564 -420 1940 -414
rect 1974 -420 1982 -334
rect 1564 -422 1982 -420
rect 1524 -436 1982 -422
rect 2030 -334 2076 1142
rect 2286 540 2724 554
rect 2286 108 2316 540
rect 2386 108 2634 540
rect 2704 108 2724 540
rect 2286 86 2724 108
rect 2942 540 3362 560
rect 2942 108 2952 540
rect 3022 108 3270 540
rect 3340 108 3362 540
rect 2942 96 3362 108
rect 2270 12 3380 24
rect 2270 -22 2282 12
rect 3374 -22 3380 12
rect 2270 -42 3380 -22
rect 2128 -312 2294 -310
rect 2030 -420 2036 -334
rect 2070 -420 2076 -334
rect 2030 -434 2076 -420
rect 2126 -334 2294 -312
rect 2126 -420 2132 -334
rect 2166 -342 2294 -334
rect 2166 -404 2246 -342
rect 2282 -390 2294 -342
rect 2282 -404 2386 -390
rect 2166 -420 2386 -404
rect 2126 -436 2386 -420
rect 1524 -437 1978 -436
rect 1524 -440 1930 -437
rect 2176 -440 2386 -436
rect 1212 -442 1335 -440
rect 1573 -442 1886 -440
rect 1212 -444 1282 -442
rect 1573 -446 1880 -442
rect 1624 -448 1880 -446
rect 1624 -450 1694 -448
rect 1959 -468 2145 -465
rect 1364 -471 1545 -469
rect 1364 -523 1370 -471
rect 1538 -523 1545 -471
rect 1364 -529 1545 -523
rect 1959 -520 1967 -468
rect 2135 -520 2145 -468
rect 1959 -527 2145 -520
rect 2228 -709 2386 -440
rect 384 -874 1566 -858
rect 384 -908 490 -874
rect 1466 -902 1566 -874
rect 2228 -860 2294 -709
rect 2228 -896 2242 -860
rect 2280 -896 2294 -860
rect 1466 -908 2012 -902
rect 2228 -906 2294 -896
rect 384 -922 2012 -908
rect 384 -936 470 -922
rect 384 -1304 406 -936
rect 440 -1304 470 -936
rect 384 -1320 470 -1304
rect 1510 -924 2012 -922
rect 1510 -936 1968 -924
rect 1510 -1304 1516 -936
rect 1550 -972 1968 -936
rect 1550 -1273 1693 -972
rect 1808 -1273 1968 -972
rect 1550 -1292 1968 -1273
rect 2002 -1292 2012 -924
rect 1550 -1304 2012 -1292
rect 1510 -1326 2012 -1304
rect 2436 -1320 2714 -1312
rect 884 -1332 1132 -1326
rect 884 -1366 934 -1332
rect 1070 -1366 1132 -1332
rect 884 -1402 1132 -1366
rect 2436 -1354 2494 -1320
rect 2626 -1354 2714 -1320
rect 222 -1404 1668 -1402
rect 2436 -1404 2714 -1354
rect 3146 -1402 3228 -42
rect 3030 -1404 3238 -1402
rect 222 -1434 3238 -1404
rect 222 -1446 1962 -1434
rect 222 -1480 400 -1446
rect 1556 -1468 1962 -1446
rect 3118 -1468 3238 -1434
rect 1556 -1480 3238 -1468
rect 222 -2573 3238 -1480
rect 222 -2734 306 -2573
rect 3154 -2734 3238 -2573
rect 222 -2837 3238 -2734
<< via1 >>
rect 150 2038 3286 2057
rect 150 1972 242 2038
rect 242 1972 314 2038
rect 314 2036 2458 2038
rect 314 2032 2018 2036
rect 314 1972 552 2032
rect 150 1966 552 1972
rect 552 1966 624 2032
rect 624 2026 1344 2032
rect 624 1966 868 2026
rect 150 1960 868 1966
rect 868 1960 940 2026
rect 940 1966 1344 2026
rect 1344 1966 1416 2032
rect 1416 1970 2018 2032
rect 2018 1970 2090 2036
rect 2090 1972 2458 2036
rect 2458 1972 2530 2038
rect 2530 1972 2752 2038
rect 2752 1972 2824 2038
rect 2824 1972 3054 2038
rect 3054 1972 3126 2038
rect 3126 1972 3286 2038
rect 2090 1970 3286 1972
rect 1416 1966 3286 1970
rect 940 1960 3286 1966
rect 150 1921 3286 1960
rect 1196 1197 1392 1538
rect 2056 1193 2249 1546
rect 1370 -476 1538 -471
rect 1370 -514 1377 -476
rect 1377 -514 1532 -476
rect 1532 -514 1538 -476
rect 1370 -523 1538 -514
rect 1967 -474 2135 -468
rect 1967 -510 1974 -474
rect 1974 -510 2132 -474
rect 2132 -510 2135 -474
rect 1967 -520 2135 -510
rect 1693 -1273 1808 -972
rect 306 -2734 3154 -2573
<< metal2 >>
rect 36 2842 3394 2927
rect 36 2658 115 2842
rect 3296 2658 3394 2842
rect 36 2057 3394 2658
rect 36 1921 150 2057
rect 3286 1921 3394 2057
rect 36 1870 3394 1921
rect -922 1565 1484 1626
rect -922 1208 -838 1565
rect -613 1538 1484 1565
rect -613 1208 1196 1538
rect -922 1197 1196 1208
rect 1392 1197 1484 1538
rect -922 1137 1484 1197
rect 1992 1546 4464 1615
rect 1992 1193 2056 1546
rect 2249 1531 4464 1546
rect 2249 1193 4154 1531
rect 1992 1174 4154 1193
rect 4379 1174 4464 1531
rect 1992 1125 4464 1174
rect -1024 -448 -731 -375
rect -812 -467 -731 -448
rect 4118 -448 4411 -375
rect -812 -471 1549 -467
rect -812 -523 1370 -471
rect 1538 -523 1549 -471
rect -812 -527 1549 -523
rect 1952 -468 4118 -462
rect 1952 -520 1967 -468
rect 2135 -520 4118 -468
rect -812 -648 -731 -527
rect 1952 -554 4118 -520
rect -1024 -709 -731 -648
rect 4330 -648 4411 -448
rect 4118 -709 4411 -648
rect 1632 -972 1891 -892
rect 1632 -1273 1693 -972
rect 1808 -1273 1891 -972
rect 1632 -1636 1891 -1273
rect 1632 -1728 4391 -1636
rect 1632 -1916 4073 -1728
rect 4287 -1916 4391 -1728
rect 1632 -1999 4391 -1916
rect 151 -2573 3297 -2515
rect 151 -2659 306 -2573
rect 151 -2825 300 -2659
rect 3154 -2734 3297 -2573
rect 3142 -2825 3297 -2734
rect 151 -2900 3297 -2825
<< via2 >>
rect 115 2658 3296 2842
rect -838 1208 -613 1565
rect 4154 1174 4379 1531
rect -1024 -648 -812 -448
rect 4118 -648 4330 -448
rect 4073 -1916 4287 -1728
rect 300 -2734 306 -2659
rect 306 -2734 3142 -2659
rect 300 -2825 3142 -2734
<< metal3 >>
rect 36 3051 3394 3193
rect 36 2853 114 3051
rect 3298 2853 3394 3051
rect 36 2842 3394 2853
rect 36 2658 115 2842
rect 3296 2658 3394 2842
rect 36 2592 3394 2658
rect -1334 1618 -555 1768
rect -1334 1162 -1213 1618
rect -740 1565 -555 1618
rect -613 1208 -555 1565
rect -740 1162 -555 1208
rect -1334 1000 -555 1162
rect 4073 1578 4681 1711
rect 4073 1531 4200 1578
rect 4073 1174 4154 1531
rect 4073 1139 4200 1174
rect 4559 1139 4681 1578
rect 4073 1006 4681 1139
rect -1059 -428 -618 -341
rect -1059 -448 -969 -428
rect -1059 -648 -1024 -448
rect -1059 -674 -969 -648
rect -699 -674 -618 -428
rect -1059 -750 -618 -674
rect 4083 -428 4524 -341
rect 4083 -448 4173 -428
rect 4083 -648 4118 -448
rect 4083 -674 4173 -648
rect 4443 -674 4524 -428
rect 4083 -750 4524 -674
rect 4003 -1682 4406 -1618
rect 4003 -1963 4061 -1682
rect 4354 -1963 4406 -1682
rect 4003 -2015 4406 -1963
rect 93 -2613 3309 -2475
rect 93 -2854 220 -2613
rect 3177 -2854 3309 -2613
rect 93 -2958 3309 -2854
<< via3 >>
rect 114 2853 3298 3051
rect -1213 1565 -740 1618
rect -1213 1208 -838 1565
rect -838 1208 -740 1565
rect -1213 1162 -740 1208
rect 4200 1531 4559 1578
rect 4200 1174 4379 1531
rect 4379 1174 4559 1531
rect 4200 1139 4559 1174
rect -969 -448 -699 -428
rect -969 -648 -812 -448
rect -812 -648 -699 -448
rect -969 -674 -699 -648
rect 4173 -448 4443 -428
rect 4173 -648 4330 -448
rect 4330 -648 4443 -448
rect 4173 -674 4443 -648
rect 4061 -1728 4354 -1682
rect 4061 -1916 4073 -1728
rect 4073 -1916 4287 -1728
rect 4287 -1916 4354 -1728
rect 4061 -1963 4354 -1916
rect 220 -2659 3177 -2613
rect 220 -2825 300 -2659
rect 300 -2825 3142 -2659
rect 3142 -2825 3177 -2659
rect 220 -2854 3177 -2825
<< metal4 >>
rect 36 3648 3405 3794
rect 36 3299 251 3648
rect 3187 3299 3405 3648
rect 36 3051 3405 3299
rect 36 2853 114 3051
rect 3298 2853 3405 3051
rect 36 2750 3405 2853
rect -1611 1785 -555 1941
rect -1611 960 -1484 1785
rect -705 960 -555 1785
rect 4033 1752 4785 1804
rect 4033 971 4095 1752
rect -1611 804 -555 960
rect -1073 -393 -598 -321
rect -1073 -718 -1021 -393
rect -665 -718 -598 -393
rect -1073 -761 -598 -718
rect 4069 -393 4544 -321
rect 4069 -718 4121 -393
rect 4477 -718 4544 -393
rect 4069 -761 4544 -718
rect 3977 -1656 4475 -1589
rect 3977 -1974 4029 -1656
rect 4417 -1974 4475 -1656
rect 3977 -2041 4475 -1974
rect 42 -2492 3389 -2395
rect 42 -2986 168 -2492
rect 3269 -2986 3389 -2492
rect 42 -3090 3389 -2986
<< via4 >>
rect 251 3299 3187 3648
rect -1484 1618 -705 1785
rect -1484 1162 -1213 1618
rect -1213 1162 -740 1618
rect -740 1162 -705 1618
rect -1484 960 -705 1162
rect 4095 1578 5000 1752
rect 4095 1139 4200 1578
rect 4200 1139 4559 1578
rect 4559 1139 5000 1578
rect 4095 697 5000 1139
rect -1021 -428 -665 -393
rect -1021 -674 -969 -428
rect -969 -674 -699 -428
rect -699 -674 -665 -428
rect -1021 -718 -665 -674
rect 4121 -428 4477 -393
rect 4121 -674 4173 -428
rect 4173 -674 4443 -428
rect 4443 -674 4477 -428
rect 4121 -718 4477 -674
rect 4029 -1682 4417 -1656
rect 4029 -1963 4061 -1682
rect 4061 -1963 4354 -1682
rect 4354 -1963 4417 -1682
rect 4029 -1974 4417 -1963
rect 168 -2613 3269 -2492
rect 168 -2854 220 -2613
rect 220 -2854 3177 -2613
rect 3177 -2854 3269 -2613
rect 168 -2986 3269 -2854
<< metal5 >>
rect -220 3648 3674 4095
rect -220 3299 251 3648
rect 3187 3299 3674 3648
rect -220 2777 3674 3299
rect -1992 1785 -532 2143
rect -1992 960 -1484 1785
rect -705 960 -532 1785
rect -1992 556 -532 960
rect 3968 1752 5464 2135
rect 3968 697 4095 1752
rect 5000 697 5464 1752
rect 3968 419 5464 697
rect -1122 -393 -508 -257
rect -1122 -718 -1021 -393
rect -665 -718 -508 -393
rect -1122 -819 -508 -718
rect 4020 -393 4634 -257
rect 4020 -718 4121 -393
rect 4477 -718 4634 -393
rect 4020 -819 4634 -718
rect 3922 -1656 4565 -1505
rect 3922 -1974 4029 -1656
rect 4417 -1974 4565 -1656
rect 3922 -2087 4565 -1974
rect -136 -2492 3561 -2263
rect -136 -2986 168 -2492
rect 3269 -2986 3561 -2492
rect -136 -3503 3561 -2986
use sky130_fd_pr__res_xhigh_po_0p35_RRCNTY  sky130_fd_pr__res_xhigh_po_0p35_RRCNTY_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606013492
transform 1 0 625 0 1 855
box -678 -908 678 908
use sky130_fd_pr__res_xhigh_po_0p35_RRCNTY  sky130_fd_pr__res_xhigh_po_0p35_RRCNTY_1
timestamp 1606013492
transform 1 0 2828 0 1 850
box -678 -908 678 908
use sky130_fd_pr__nfet_01v8_lvt_PZT9H9  sky130_fd_pr__nfet_01v8_lvt_PZT9H9_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606079819
transform 1 0 2051 0 1 -371
box -263 -265 263 265
use sky130_fd_pr__nfet_01v8_lvt_PZT9H9  sky130_fd_pr__nfet_01v8_lvt_PZT9H9_1
timestamp 1606079819
transform 1 0 1453 0 1 -377
box -263 -265 263 265
use sky130_fd_pr__nfet_01v8_lvt_F9NR5A  sky130_fd_pr__nfet_01v8_lvt_F9NR5A_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606079819
transform 0 1 2542 -1 0 -1106
box -396 -710 396 710
use sky130_fd_pr__nfet_01v8_lvt_F9NR5A  sky130_fd_pr__nfet_01v8_lvt_F9NR5A_1
timestamp 1606079819
transform 0 1 976 -1 0 -1120
box -396 -710 396 710
<< labels >>
rlabel via1 1676 1966 1770 2038 1 Vdd
port 1 n
rlabel metal1 2018 1326 2108 1452 1 ON2a
port 2 n
rlabel metal1 1370 1334 1460 1460 1 ON1a
port 3 n
rlabel poly 1996 -272 2014 -248 1 VN
port 5 n
rlabel metal1 1720 -1526 1794 -1482 1 Gnd
port 6 n
rlabel via1 1720 -1144 1792 -1080 1 vbiasn
port 7 n
rlabel metal1 2244 -690 2270 -666 1 Itail_a
rlabel poly 1390 -276 1408 -252 1 VP
port 4 n
<< end >>
