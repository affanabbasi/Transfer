magic
tech sky130A
magscale 1 2
timestamp 1606812005
<< metal1 >>
rect 226738 -32043 357511 -31948
rect 226738 -32400 354392 -32043
rect 357432 -32400 357511 -32043
rect 226738 -32479 357511 -32400
rect 320307 -32733 322284 -32479
rect 234229 -43727 286945 -40124
rect 234229 -45211 234764 -43727
rect 286475 -45211 286945 -43727
rect 234229 -45806 286945 -45211
<< via1 >>
rect 354392 -32400 357432 -32043
rect 236556 -39428 236637 -39363
rect 234764 -45211 286475 -43727
<< metal2 >>
rect 54068 382528 95797 384682
rect 54068 375428 55689 382528
rect 54068 374841 58946 375428
rect 63466 374856 64082 375443
rect 73283 375165 74904 382528
rect 94176 376752 95797 382528
rect 94176 376165 99689 376752
rect 73283 374578 78161 375165
rect 5151 369751 6242 373268
rect 63369 369751 64414 374079
rect 77713 369751 78139 374217
rect 5151 368243 78139 369751
rect -19560 -21048 173239 -20510
rect -19560 -29114 -19099 -21048
rect -11205 -29114 173239 -21048
rect -19560 -29621 173239 -29114
rect 354300 -32043 357511 -31920
rect 354300 -32400 354392 -32043
rect 357432 -32400 357511 -32043
rect 354300 -33958 357511 -32400
rect 234261 -39363 236666 -38413
rect 234261 -39428 236556 -39363
rect 236637 -39428 236666 -39363
rect 234261 -39463 236666 -39428
rect 234229 -43637 286945 -43222
rect 234229 -45351 234646 -43637
rect 286559 -45351 286945 -43637
rect 234229 -45806 286945 -45351
<< via2 >>
rect -19099 -29114 -11205 -21048
rect 234646 -43727 286559 -43637
rect 234646 -45211 234764 -43727
rect 234764 -45211 286475 -43727
rect 286475 -45211 286559 -43727
rect 234646 -45351 286559 -45211
<< metal3 >>
rect -19560 380290 38105 381411
rect -19560 -21048 -10715 380290
rect -3560 378399 -2469 380290
rect 37014 378002 38105 380290
rect 67277 381251 91037 383003
rect 67277 375443 68898 381251
rect 63466 374856 68898 375443
rect 89478 375901 91037 381251
rect 100799 375901 101451 376667
rect 89478 375314 101451 375901
rect 89478 375217 91037 375314
rect 83993 374610 91037 375217
rect -19560 -29114 -19099 -21048
rect -11205 -29114 -10715 -21048
rect -19560 -29621 -10715 -29114
rect 234229 -43530 286945 -43222
rect 234229 -45474 234540 -43530
rect 286648 -45474 286945 -43530
rect 234229 -45806 286945 -45474
<< via3 >>
rect 234540 -43637 286648 -43530
rect 234540 -45351 234646 -43637
rect 234646 -45351 286559 -43637
rect 286559 -45351 286648 -43637
rect 234540 -45474 286648 -45351
<< metal4 >>
rect 95894 360081 97123 373638
rect -34915 349108 97123 360081
rect -34915 -51999 -25820 349108
rect 185527 -36496 196607 -33773
rect 192914 -51999 196607 -36496
rect 234229 -43417 286945 -43222
rect 234229 -45623 234401 -43417
rect 286756 -45623 286945 -43417
rect 234229 -45806 286945 -45623
rect -34915 -57298 196607 -51999
<< via4 >>
rect 234401 -43530 286756 -43417
rect 234401 -45474 234540 -43530
rect 234540 -45474 286648 -43530
rect 286648 -45474 286756 -43530
rect 234401 -45623 286756 -45474
<< metal5 >>
rect 14438 385214 112146 389734
rect 14438 377432 16116 385214
rect 39590 378351 40052 385214
rect 59233 379762 63127 385214
rect 80138 380492 82041 385214
rect 96486 381115 97126 385214
rect 14470 364767 15874 374282
rect 39447 364767 40212 373690
rect 59219 364767 63111 372295
rect 80247 364767 82311 372084
rect 97955 364767 98612 372645
rect -52977 360247 112178 364767
rect -52977 -43222 -47130 360247
rect 178831 -29552 354135 -24375
rect 238719 -31764 239616 -29552
rect 317049 -34344 317515 -29552
rect 353386 -34766 354135 -29552
rect 184807 -43222 187145 -38239
rect 317046 -43222 317512 -37088
rect 354350 -43222 357843 -36038
rect -52977 -43417 358077 -43222
rect -52977 -45623 234401 -43417
rect 286756 -45623 358077 -43417
rect -52977 -46201 358077 -45623
use RO  RO_0 ~/CustomFlow/magic/Work-main/layouts/RingOscillator
timestamp 1606670916
transform 1 0 354350 0 1 -35359
box -918 -687 4384 1644
use BiasVCO  BiasVCO_0 ~/CustomFlow/magic/Work-main/layouts/VCO/BiasVCO
timestamp 1606672880
transform 1 0 317789 0 1 -35727
box -743 -1581 14424 3042
use Delay_Top  Delay_Top_0
timestamp 1606686671
transform 1 0 223681 0 1 -40002
box 3057 -128 65878 14314
use PA_1  PA_1_0
timestamp 1606531739
transform 1 0 15084 0 1 -7863
box 0 -31847 352952 379374
use LVDStop  LVDStop_0 ~/CustomFlow/magic/Work-main/layouts/LVDS/lvdstop
timestamp 1606674334
transform 1 0 -2045 0 1 373048
box -1515 0 20087 5918
use LVDSBias_Top  LVDSBias_Top_0
timestamp 1606670916
transform 1 0 39318 0 1 377835
box -3702 -5224 3568 842
use LVDS1_Top  LVDS1_Top_0
timestamp 1606621314
transform 1 0 59453 0 1 375677
box -1992 -3503 5464 4095
use LVDS2_Top  LVDS2_Top_0
timestamp 1606674334
transform 1 0 78399 0 1 375538
box -694 -3510 6019 4973
use foldedcascode1  foldedcascode1_0
timestamp 1606790247
transform 1 0 100046 0 1 376620
box -3600 -4460 11100 4600
<< labels >>
rlabel metal5 350574 -28978 353470 -25117 1 p_vgate
port 1 n
rlabel space 355778 341564 365860 351484 1 pa_vdd
port 2 n
rlabel metal5 15373 386177 18490 389054 1 p_vdd
port 3 n
rlabel metal5 354549 -46011 357666 -43134 1 p_vss
port 4 n
rlabel metal4 -33179 350269 -26691 358785 1 p_isrc
port 5 n
rlabel space 358217 -35355 358690 -34477 1 ro_out
port 6 n
rlabel space 320328 -37256 320662 -36917 1 selfb_vinit
port 7 n
rlabel space 317084 -36228 317493 -35818 1 selfb_vbn
port 8 n
rlabel space 317085 -35318 317474 -34934 1 inv1in
port 9 n
rlabel space 232970 -35488 233359 -35104 1 dvco_outn
port 10 n
rlabel space 229038 -36503 229427 -36119 1 dvco_outp
port 11 n
rlabel metal2 234466 -39151 234911 -38685 1 dvco_vbn
port 12 n
rlabel space 183113 -31067 183558 -30601 1 pa_rnode
port 13 n
rlabel space 164633 -17763 168822 -12003 1 pa_out
port 14 n
rlabel space 17146 375540 17814 376244 1 lvdstop_out
port 15 n
rlabel space -3189 376859 -2851 377183 1 lvdstop_inp
port 16 n
rlabel space -3154 375288 -2816 375612 1 lvdstop_inn
port 17 n
rlabel metal2 5345 368405 6973 369580 1 lvds_vbiasn
port 18 n
rlabel space 35734 376337 35891 376501 1 lvdsbias_inp
port 19 n
rlabel space 35734 374811 35891 374975 1 lvdsbias_inn
port 20 n
rlabel space 42549 376929 42755 377132 1 lvdsbias_vp
port 21 n
rlabel space 42549 375903 42755 376106 1 lvdsbias_vn
port 22 n
rlabel space 57700 376413 58664 377615 1 lvds1_on1a
port 23 n
rlabel space 63680 376312 64644 377514 1 lvds1_on2a
port 24 n
rlabel metal2 54419 382763 57012 384413 1 lvds_vp
port 25 n
rlabel metal3 67486 381298 70113 382427 1 lvds_vn
port 26 n
rlabel space 77777 375393 78027 375661 1 lvds2_on2b
port 27 n
rlabel space 84072 375393 84322 375661 1 lvds2_on1b
port 28 n
rlabel space 108574 377846 109032 378241 1 fc_out
port 29 n
rlabel metal2 354618 -33602 357246 -32661 1 ocs_vdd
port 30 n
<< end >>
