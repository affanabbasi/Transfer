magic
tech sky130A
timestamp 1606452767
<< metal4 >>
rect -136800 -5800 -119100 89100
rect -136800 -13200 -136500 -5800
rect -119400 -13200 -119100 -5800
rect -136800 -13500 -119100 -13200
<< via4 >>
rect -136500 -13200 -119400 -5800
<< metal5 >>
rect -216300 73500 -39900 81500
rect -216300 -59500 -208300 73500
rect -198300 55500 -57900 63500
rect -198300 -41500 -190300 55500
rect -180300 37500 -75900 45500
rect -180300 -23500 -172300 37500
rect -162300 19500 -93900 27500
rect -162300 -5500 -154300 19500
rect -162300 -5800 -119100 -5500
rect -162300 -13200 -136500 -5800
rect -119400 -13200 -119100 -5800
rect -162300 -13500 -119100 -13200
rect -101900 -23500 -93900 19500
rect -180300 -31500 -93900 -23500
rect -83900 -41500 -75900 37500
rect -198300 -49500 -75900 -41500
rect -65900 -59500 -57900 55500
rect -216300 -67500 -57900 -59500
rect -47900 -77500 -39900 73500
rect -141400 -85500 -39900 -77500
<< end >>
