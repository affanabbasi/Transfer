magic
tech sky130A
timestamp 1606578544
<< pwell >>
rect -885 -455 885 455
<< nmos >>
rect -787 -350 -587 350
rect -558 -350 -358 350
rect -329 -350 -129 350
rect -100 -350 100 350
rect 129 -350 329 350
rect 358 -350 558 350
rect 587 -350 787 350
<< ndiff >>
rect -816 344 -787 350
rect -816 -344 -810 344
rect -793 -344 -787 344
rect -816 -350 -787 -344
rect -587 344 -558 350
rect -587 -344 -581 344
rect -564 -344 -558 344
rect -587 -350 -558 -344
rect -358 344 -329 350
rect -358 -344 -352 344
rect -335 -344 -329 344
rect -358 -350 -329 -344
rect -129 344 -100 350
rect -129 -344 -123 344
rect -106 -344 -100 344
rect -129 -350 -100 -344
rect 100 344 129 350
rect 100 -344 106 344
rect 123 -344 129 344
rect 100 -350 129 -344
rect 329 344 358 350
rect 329 -344 335 344
rect 352 -344 358 344
rect 329 -350 358 -344
rect 558 344 587 350
rect 558 -344 564 344
rect 581 -344 587 344
rect 558 -350 587 -344
rect 787 344 816 350
rect 787 -344 793 344
rect 810 -344 816 344
rect 787 -350 816 -344
<< ndiffc >>
rect -810 -344 -793 344
rect -581 -344 -564 344
rect -352 -344 -335 344
rect -123 -344 -106 344
rect 106 -344 123 344
rect 335 -344 352 344
rect 564 -344 581 344
rect 793 -344 810 344
<< psubdiff >>
rect -867 420 -819 437
rect 819 420 867 437
rect -867 389 -850 420
rect 850 389 867 420
rect -867 -420 -850 -389
rect 850 -420 867 -389
rect -867 -437 -819 -420
rect 819 -437 867 -420
<< psubdiffcont >>
rect -819 420 819 437
rect -867 -389 -850 389
rect 850 -389 867 389
rect -819 -437 819 -420
<< poly >>
rect -787 386 -587 394
rect -787 369 -779 386
rect -595 369 -587 386
rect -787 350 -587 369
rect -558 386 -358 394
rect -558 369 -550 386
rect -366 369 -358 386
rect -558 350 -358 369
rect -329 386 -129 394
rect -329 369 -321 386
rect -137 369 -129 386
rect -329 350 -129 369
rect -100 386 100 394
rect -100 369 -92 386
rect 92 369 100 386
rect -100 350 100 369
rect 129 386 329 394
rect 129 369 137 386
rect 321 369 329 386
rect 129 350 329 369
rect 358 386 558 394
rect 358 369 366 386
rect 550 369 558 386
rect 358 350 558 369
rect 587 386 787 394
rect 587 369 595 386
rect 779 369 787 386
rect 587 350 787 369
rect -787 -369 -587 -350
rect -787 -386 -779 -369
rect -595 -386 -587 -369
rect -787 -394 -587 -386
rect -558 -369 -358 -350
rect -558 -386 -550 -369
rect -366 -386 -358 -369
rect -558 -394 -358 -386
rect -329 -369 -129 -350
rect -329 -386 -321 -369
rect -137 -386 -129 -369
rect -329 -394 -129 -386
rect -100 -369 100 -350
rect -100 -386 -92 -369
rect 92 -386 100 -369
rect -100 -394 100 -386
rect 129 -369 329 -350
rect 129 -386 137 -369
rect 321 -386 329 -369
rect 129 -394 329 -386
rect 358 -369 558 -350
rect 358 -386 366 -369
rect 550 -386 558 -369
rect 358 -394 558 -386
rect 587 -369 787 -350
rect 587 -386 595 -369
rect 779 -386 787 -369
rect 587 -394 787 -386
<< polycont >>
rect -779 369 -595 386
rect -550 369 -366 386
rect -321 369 -137 386
rect -92 369 92 386
rect 137 369 321 386
rect 366 369 550 386
rect 595 369 779 386
rect -779 -386 -595 -369
rect -550 -386 -366 -369
rect -321 -386 -137 -369
rect -92 -386 92 -369
rect 137 -386 321 -369
rect 366 -386 550 -369
rect 595 -386 779 -369
<< locali >>
rect -867 420 -819 437
rect 819 420 867 437
rect -867 389 -850 420
rect 850 389 867 420
rect -787 369 -779 386
rect -595 369 -587 386
rect -558 369 -550 386
rect -366 369 -358 386
rect -329 369 -321 386
rect -137 369 -129 386
rect -100 369 -92 386
rect 92 369 100 386
rect 129 369 137 386
rect 321 369 329 386
rect 358 369 366 386
rect 550 369 558 386
rect 587 369 595 386
rect 779 369 787 386
rect -810 344 -793 352
rect -810 -352 -793 -344
rect -581 344 -564 352
rect -581 -352 -564 -344
rect -352 344 -335 352
rect -352 -352 -335 -344
rect -123 344 -106 352
rect -123 -352 -106 -344
rect 106 344 123 352
rect 106 -352 123 -344
rect 335 344 352 352
rect 335 -352 352 -344
rect 564 344 581 352
rect 564 -352 581 -344
rect 793 344 810 352
rect 793 -352 810 -344
rect -787 -386 -779 -369
rect -595 -386 -587 -369
rect -558 -386 -550 -369
rect -366 -386 -358 -369
rect -329 -386 -321 -369
rect -137 -386 -129 -369
rect -100 -386 -92 -369
rect 92 -386 100 -369
rect 129 -386 137 -369
rect 321 -386 329 -369
rect 358 -386 366 -369
rect 550 -386 558 -369
rect 587 -386 595 -369
rect 779 -386 787 -369
rect -867 -420 -850 -389
rect 850 -420 867 -389
rect -867 -437 -819 -420
rect 819 -437 867 -420
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -858 -428 858 428
string parameters w 7 l 2 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
