magic
tech sky130A
magscale 1 2
timestamp 1606422944
<< pwell >>
rect 35469 1159 35503 3135
<< ndiff >>
rect 35469 1159 35503 3135
<< locali >>
rect 29165 3186 29170 3219
rect 38624 3186 38639 3219
rect 29165 3185 38639 3186
rect 29069 1102 38543 1109
rect 29069 1075 29070 1102
rect 38524 1075 38543 1102
<< viali >>
rect 29170 3186 38624 3226
rect 29037 1159 29071 3135
rect 29133 1159 29167 3135
rect 29229 1159 29263 3135
rect 29325 1159 29359 3135
rect 29421 1159 29455 3135
rect 29517 1159 29551 3135
rect 29613 1159 29647 3135
rect 29709 1159 29743 3135
rect 29805 1159 29839 3135
rect 29901 1159 29935 3135
rect 29997 1159 30031 3135
rect 30093 1159 30127 3135
rect 30189 1159 30223 3135
rect 30285 1159 30319 3135
rect 30381 1159 30415 3135
rect 30477 1159 30511 3135
rect 30573 1159 30607 3135
rect 30669 1159 30703 3135
rect 30765 1159 30799 3135
rect 30861 1159 30895 3135
rect 30957 1159 30991 3135
rect 31053 1159 31087 3135
rect 31149 1159 31183 3135
rect 31245 1159 31279 3135
rect 31341 1159 31375 3135
rect 31437 1159 31471 3135
rect 31533 1159 31567 3135
rect 31629 1159 31663 3135
rect 31725 1159 31759 3135
rect 31821 1159 31855 3135
rect 31917 1159 31951 3135
rect 32013 1159 32047 3135
rect 32109 1159 32143 3135
rect 32205 1159 32239 3135
rect 32301 1159 32335 3135
rect 32397 1159 32431 3135
rect 32493 1159 32527 3135
rect 32589 1159 32623 3135
rect 32685 1159 32719 3135
rect 32781 1159 32815 3135
rect 32877 1159 32911 3135
rect 32973 1159 33007 3135
rect 33069 1159 33103 3135
rect 33165 1159 33199 3135
rect 33261 1159 33295 3135
rect 33357 1159 33391 3135
rect 33453 1159 33487 3135
rect 33549 1159 33583 3135
rect 33645 1159 33679 3135
rect 33741 1159 33775 3135
rect 33837 1159 33871 3135
rect 33933 1159 33967 3135
rect 34029 1159 34063 3135
rect 34125 1159 34159 3135
rect 34221 1159 34255 3135
rect 34317 1159 34351 3135
rect 34413 1159 34447 3135
rect 34509 1159 34543 3135
rect 34605 1159 34639 3135
rect 34701 1159 34735 3135
rect 34797 1159 34831 3135
rect 34893 1159 34927 3135
rect 34989 1159 35023 3135
rect 35085 1159 35119 3135
rect 35181 1159 35215 3135
rect 35277 1159 35311 3135
rect 35373 1159 35407 3135
rect 35469 1159 35503 3135
rect 35565 1159 35599 3135
rect 35661 1159 35695 3135
rect 35757 1159 35791 3135
rect 35853 1159 35887 3135
rect 35949 1159 35983 3135
rect 36045 1159 36079 3135
rect 36141 1159 36175 3135
rect 36237 1159 36271 3135
rect 36333 1159 36367 3135
rect 36429 1159 36463 3135
rect 36525 1159 36559 3135
rect 36621 1159 36655 3135
rect 36717 1159 36751 3135
rect 36813 1159 36847 3135
rect 36909 1159 36943 3135
rect 37005 1159 37039 3135
rect 37101 1159 37135 3135
rect 37197 1159 37231 3135
rect 37293 1159 37327 3135
rect 37389 1159 37423 3135
rect 37485 1159 37519 3135
rect 37581 1159 37615 3135
rect 37677 1159 37711 3135
rect 37773 1159 37807 3135
rect 37869 1159 37903 3135
rect 37965 1159 37999 3135
rect 38061 1159 38095 3135
rect 38157 1159 38191 3135
rect 38253 1159 38287 3135
rect 38349 1159 38383 3135
rect 38445 1159 38479 3135
rect 38541 1159 38575 3135
rect 38637 1158 38671 3134
rect 29070 1062 38524 1102
<< metal1 >>
rect 29140 3226 38986 3250
rect 29140 3186 29170 3226
rect 38624 3186 38986 3226
rect 29140 3180 38986 3186
rect 29140 3176 29186 3180
rect 29025 3135 29083 3147
rect 29025 1159 29028 3135
rect 29080 1159 29083 3135
rect 29025 1147 29083 1159
rect 29121 3135 29179 3147
rect 29121 1159 29124 3135
rect 29176 1159 29179 3135
rect 29121 1147 29179 1159
rect 29217 3135 29275 3147
rect 29217 1159 29220 3135
rect 29272 1159 29275 3135
rect 29217 1147 29275 1159
rect 29316 3135 29368 3147
rect 29316 1147 29368 1159
rect 29409 3135 29467 3147
rect 29409 1159 29412 3135
rect 29464 1159 29467 3135
rect 29409 1147 29467 1159
rect 29505 3135 29563 3147
rect 29505 1159 29508 3135
rect 29560 1159 29563 3135
rect 29505 1147 29563 1159
rect 29601 3135 29659 3147
rect 29601 1159 29604 3135
rect 29656 1159 29659 3135
rect 29601 1147 29659 1159
rect 29700 3135 29752 3147
rect 29700 1147 29752 1159
rect 29793 3135 29851 3147
rect 29793 1159 29796 3135
rect 29848 1159 29851 3135
rect 29793 1147 29851 1159
rect 29889 3135 29947 3147
rect 29889 1159 29892 3135
rect 29944 1159 29947 3135
rect 29889 1147 29947 1159
rect 29985 3135 30043 3147
rect 29985 1159 29988 3135
rect 30040 1159 30043 3135
rect 29985 1147 30043 1159
rect 30084 3135 30136 3147
rect 30084 1147 30136 1159
rect 30177 3135 30235 3147
rect 30177 1159 30180 3135
rect 30232 1159 30235 3135
rect 30177 1147 30235 1159
rect 30273 3135 30331 3147
rect 30273 1159 30276 3135
rect 30328 1159 30331 3135
rect 30273 1147 30331 1159
rect 30369 3135 30427 3147
rect 30369 1159 30372 3135
rect 30424 1159 30427 3135
rect 30369 1147 30427 1159
rect 30468 3135 30520 3147
rect 30468 1147 30520 1159
rect 30561 3135 30619 3147
rect 30561 1159 30564 3135
rect 30616 1159 30619 3135
rect 30561 1147 30619 1159
rect 30657 3135 30715 3147
rect 30657 1159 30660 3135
rect 30712 1159 30715 3135
rect 30657 1147 30715 1159
rect 30753 3135 30811 3147
rect 30753 1159 30756 3135
rect 30808 1159 30811 3135
rect 30753 1147 30811 1159
rect 30852 3135 30904 3147
rect 30852 1147 30904 1159
rect 30945 3135 31003 3147
rect 30945 1159 30948 3135
rect 31000 1159 31003 3135
rect 30945 1147 31003 1159
rect 31041 3135 31099 3147
rect 31041 1159 31044 3135
rect 31096 1159 31099 3135
rect 31041 1147 31099 1159
rect 31137 3135 31195 3147
rect 31137 1159 31140 3135
rect 31192 1159 31195 3135
rect 31137 1147 31195 1159
rect 31236 3135 31288 3147
rect 31236 1147 31288 1159
rect 31329 3135 31387 3147
rect 31329 1159 31332 3135
rect 31384 1159 31387 3135
rect 31329 1147 31387 1159
rect 31425 3135 31483 3147
rect 31425 1159 31428 3135
rect 31480 1159 31483 3135
rect 31425 1147 31483 1159
rect 31521 3135 31579 3147
rect 31521 1159 31524 3135
rect 31576 1159 31579 3135
rect 31521 1147 31579 1159
rect 31620 3135 31672 3147
rect 31620 1147 31672 1159
rect 31713 3135 31771 3147
rect 31713 1159 31716 3135
rect 31768 1159 31771 3135
rect 31713 1147 31771 1159
rect 31809 3135 31867 3147
rect 31809 1159 31812 3135
rect 31864 1159 31867 3135
rect 31809 1147 31867 1159
rect 31905 3135 31963 3147
rect 31905 1159 31908 3135
rect 31960 1159 31963 3135
rect 31905 1147 31963 1159
rect 32004 3135 32056 3147
rect 32004 1147 32056 1159
rect 32097 3135 32155 3147
rect 32097 1159 32100 3135
rect 32152 1159 32155 3135
rect 32097 1147 32155 1159
rect 32193 3135 32251 3147
rect 32193 1159 32196 3135
rect 32248 1159 32251 3135
rect 32193 1147 32251 1159
rect 32289 3135 32347 3147
rect 32289 1159 32292 3135
rect 32344 1159 32347 3135
rect 32289 1147 32347 1159
rect 32388 3135 32440 3147
rect 32388 1147 32440 1159
rect 32481 3135 32539 3147
rect 32481 1159 32484 3135
rect 32536 1159 32539 3135
rect 32481 1147 32539 1159
rect 32577 3135 32635 3147
rect 32577 1159 32580 3135
rect 32632 1159 32635 3135
rect 32577 1147 32635 1159
rect 32673 3135 32731 3147
rect 32673 1159 32676 3135
rect 32728 1159 32731 3135
rect 32673 1147 32731 1159
rect 32772 3135 32824 3147
rect 32772 1147 32824 1159
rect 32865 3135 32923 3147
rect 32865 1159 32868 3135
rect 32920 1159 32923 3135
rect 32865 1147 32923 1159
rect 32961 3135 33019 3147
rect 32961 1159 32964 3135
rect 33016 1159 33019 3135
rect 32961 1147 33019 1159
rect 33057 3135 33115 3147
rect 33057 1159 33060 3135
rect 33112 1159 33115 3135
rect 33057 1147 33115 1159
rect 33156 3135 33208 3147
rect 33156 1147 33208 1159
rect 33249 3135 33307 3147
rect 33249 1159 33252 3135
rect 33304 1159 33307 3135
rect 33249 1147 33307 1159
rect 33345 3135 33403 3147
rect 33345 1159 33348 3135
rect 33400 1159 33403 3135
rect 33345 1147 33403 1159
rect 33441 3135 33499 3147
rect 33441 1159 33444 3135
rect 33496 1159 33499 3135
rect 33441 1147 33499 1159
rect 33540 3135 33592 3147
rect 33540 1147 33592 1159
rect 33633 3135 33691 3147
rect 33633 1159 33636 3135
rect 33688 1159 33691 3135
rect 33633 1147 33691 1159
rect 33729 3135 33787 3147
rect 33729 1159 33732 3135
rect 33784 1159 33787 3135
rect 33729 1147 33787 1159
rect 33825 3135 33883 3147
rect 33825 1159 33828 3135
rect 33880 1159 33883 3135
rect 33825 1147 33883 1159
rect 33924 3135 33976 3147
rect 33924 1147 33976 1159
rect 34017 3135 34075 3147
rect 34017 1159 34020 3135
rect 34072 1159 34075 3135
rect 34017 1147 34075 1159
rect 34113 3135 34171 3147
rect 34113 1159 34116 3135
rect 34168 1159 34171 3135
rect 34113 1147 34171 1159
rect 34209 3135 34267 3147
rect 34209 1159 34212 3135
rect 34264 1159 34267 3135
rect 34209 1147 34267 1159
rect 34308 3135 34360 3147
rect 34308 1147 34360 1159
rect 34401 3135 34459 3147
rect 34401 1159 34404 3135
rect 34456 1159 34459 3135
rect 34401 1147 34459 1159
rect 34497 3135 34555 3147
rect 34497 1159 34500 3135
rect 34552 1159 34555 3135
rect 34497 1147 34555 1159
rect 34593 3135 34651 3147
rect 34593 1159 34596 3135
rect 34648 1159 34651 3135
rect 34593 1147 34651 1159
rect 34692 3135 34744 3147
rect 34692 1147 34744 1159
rect 34785 3135 34843 3147
rect 34785 1159 34788 3135
rect 34840 1159 34843 3135
rect 34785 1147 34843 1159
rect 34881 3135 34939 3147
rect 34881 1159 34884 3135
rect 34936 1159 34939 3135
rect 34881 1147 34939 1159
rect 34977 3135 35035 3147
rect 34977 1159 34980 3135
rect 35032 1159 35035 3135
rect 34977 1147 35035 1159
rect 35076 3135 35128 3147
rect 35076 1147 35128 1159
rect 35169 3135 35227 3147
rect 35169 1159 35172 3135
rect 35224 1159 35227 3135
rect 35169 1147 35227 1159
rect 35265 3135 35323 3147
rect 35265 1159 35268 3135
rect 35320 1159 35323 3135
rect 35265 1147 35323 1159
rect 35361 3135 35419 3147
rect 35361 1159 35364 3135
rect 35416 1159 35419 3135
rect 35361 1147 35419 1159
rect 35460 3135 35512 3147
rect 35460 1147 35512 1159
rect 35553 3135 35611 3147
rect 35553 1159 35556 3135
rect 35608 1159 35611 3135
rect 35553 1147 35611 1159
rect 35649 3135 35707 3147
rect 35649 1159 35652 3135
rect 35704 1159 35707 3135
rect 35649 1147 35707 1159
rect 35745 3135 35803 3147
rect 35745 1159 35748 3135
rect 35800 1159 35803 3135
rect 35745 1147 35803 1159
rect 35844 3135 35896 3147
rect 35844 1147 35896 1159
rect 35937 3135 35995 3147
rect 35937 1159 35940 3135
rect 35992 1159 35995 3135
rect 35937 1147 35995 1159
rect 36033 3135 36091 3147
rect 36033 1159 36036 3135
rect 36088 1159 36091 3135
rect 36033 1147 36091 1159
rect 36129 3135 36187 3147
rect 36129 1159 36132 3135
rect 36184 1159 36187 3135
rect 36129 1147 36187 1159
rect 36228 3135 36280 3147
rect 36228 1147 36280 1159
rect 36321 3135 36379 3147
rect 36321 1159 36324 3135
rect 36376 1159 36379 3135
rect 36321 1147 36379 1159
rect 36417 3135 36475 3147
rect 36417 1159 36420 3135
rect 36472 1159 36475 3135
rect 36417 1147 36475 1159
rect 36513 3135 36571 3147
rect 36513 1159 36516 3135
rect 36568 1159 36571 3135
rect 36513 1147 36571 1159
rect 36612 3135 36664 3147
rect 36612 1147 36664 1159
rect 36705 3135 36763 3147
rect 36705 1159 36708 3135
rect 36760 1159 36763 3135
rect 36705 1147 36763 1159
rect 36801 3135 36859 3147
rect 36801 1159 36804 3135
rect 36856 1159 36859 3135
rect 36801 1147 36859 1159
rect 36897 3135 36955 3147
rect 36897 1159 36900 3135
rect 36952 1159 36955 3135
rect 36897 1147 36955 1159
rect 36996 3135 37048 3147
rect 36996 1147 37048 1159
rect 37089 3135 37147 3147
rect 37089 1159 37092 3135
rect 37144 1159 37147 3135
rect 37089 1147 37147 1159
rect 37185 3135 37243 3147
rect 37185 1159 37188 3135
rect 37240 1159 37243 3135
rect 37185 1147 37243 1159
rect 37281 3135 37339 3147
rect 37281 1159 37284 3135
rect 37336 1159 37339 3135
rect 37281 1147 37339 1159
rect 37380 3135 37432 3147
rect 37380 1147 37432 1159
rect 37473 3135 37531 3147
rect 37473 1159 37476 3135
rect 37528 1159 37531 3135
rect 37473 1147 37531 1159
rect 37569 3135 37627 3147
rect 37569 1159 37572 3135
rect 37624 1159 37627 3135
rect 37569 1147 37627 1159
rect 37665 3135 37723 3147
rect 37665 1159 37668 3135
rect 37720 1159 37723 3135
rect 37665 1147 37723 1159
rect 37764 3135 37816 3147
rect 37764 1147 37816 1159
rect 37857 3135 37915 3147
rect 37857 1159 37860 3135
rect 37912 1159 37915 3135
rect 37857 1147 37915 1159
rect 37953 3135 38011 3147
rect 37953 1159 37956 3135
rect 38008 1159 38011 3135
rect 37953 1147 38011 1159
rect 38049 3135 38107 3147
rect 38049 1159 38052 3135
rect 38104 1159 38107 3135
rect 38049 1147 38107 1159
rect 38148 3135 38200 3147
rect 38148 1147 38200 1159
rect 38241 3135 38299 3147
rect 38241 1159 38244 3135
rect 38296 1159 38299 3135
rect 38241 1147 38299 1159
rect 38337 3135 38395 3147
rect 38337 1159 38340 3135
rect 38392 1159 38395 3135
rect 38337 1147 38395 1159
rect 38433 3135 38491 3147
rect 38433 1159 38436 3135
rect 38488 1159 38491 3135
rect 38433 1147 38491 1159
rect 38532 3135 38584 3147
rect 38532 1147 38584 1159
rect 38625 3134 38683 3146
rect 38625 1158 38628 3134
rect 38680 1158 38683 3134
rect 38625 1146 38683 1158
rect 38912 1112 38986 3180
rect 29070 1110 38986 1112
rect 29040 1102 38986 1110
rect 29040 1062 29070 1102
rect 38524 1062 38986 1102
rect 29040 1042 38986 1062
<< via1 >>
rect 29028 1159 29037 3135
rect 29037 1159 29071 3135
rect 29071 1159 29080 3135
rect 29124 1159 29133 3135
rect 29133 1159 29167 3135
rect 29167 1159 29176 3135
rect 29220 1159 29229 3135
rect 29229 1159 29263 3135
rect 29263 1159 29272 3135
rect 29316 1159 29325 3135
rect 29325 1159 29359 3135
rect 29359 1159 29368 3135
rect 29412 1159 29421 3135
rect 29421 1159 29455 3135
rect 29455 1159 29464 3135
rect 29508 1159 29517 3135
rect 29517 1159 29551 3135
rect 29551 1159 29560 3135
rect 29604 1159 29613 3135
rect 29613 1159 29647 3135
rect 29647 1159 29656 3135
rect 29700 1159 29709 3135
rect 29709 1159 29743 3135
rect 29743 1159 29752 3135
rect 29796 1159 29805 3135
rect 29805 1159 29839 3135
rect 29839 1159 29848 3135
rect 29892 1159 29901 3135
rect 29901 1159 29935 3135
rect 29935 1159 29944 3135
rect 29988 1159 29997 3135
rect 29997 1159 30031 3135
rect 30031 1159 30040 3135
rect 30084 1159 30093 3135
rect 30093 1159 30127 3135
rect 30127 1159 30136 3135
rect 30180 1159 30189 3135
rect 30189 1159 30223 3135
rect 30223 1159 30232 3135
rect 30276 1159 30285 3135
rect 30285 1159 30319 3135
rect 30319 1159 30328 3135
rect 30372 1159 30381 3135
rect 30381 1159 30415 3135
rect 30415 1159 30424 3135
rect 30468 1159 30477 3135
rect 30477 1159 30511 3135
rect 30511 1159 30520 3135
rect 30564 1159 30573 3135
rect 30573 1159 30607 3135
rect 30607 1159 30616 3135
rect 30660 1159 30669 3135
rect 30669 1159 30703 3135
rect 30703 1159 30712 3135
rect 30756 1159 30765 3135
rect 30765 1159 30799 3135
rect 30799 1159 30808 3135
rect 30852 1159 30861 3135
rect 30861 1159 30895 3135
rect 30895 1159 30904 3135
rect 30948 1159 30957 3135
rect 30957 1159 30991 3135
rect 30991 1159 31000 3135
rect 31044 1159 31053 3135
rect 31053 1159 31087 3135
rect 31087 1159 31096 3135
rect 31140 1159 31149 3135
rect 31149 1159 31183 3135
rect 31183 1159 31192 3135
rect 31236 1159 31245 3135
rect 31245 1159 31279 3135
rect 31279 1159 31288 3135
rect 31332 1159 31341 3135
rect 31341 1159 31375 3135
rect 31375 1159 31384 3135
rect 31428 1159 31437 3135
rect 31437 1159 31471 3135
rect 31471 1159 31480 3135
rect 31524 1159 31533 3135
rect 31533 1159 31567 3135
rect 31567 1159 31576 3135
rect 31620 1159 31629 3135
rect 31629 1159 31663 3135
rect 31663 1159 31672 3135
rect 31716 1159 31725 3135
rect 31725 1159 31759 3135
rect 31759 1159 31768 3135
rect 31812 1159 31821 3135
rect 31821 1159 31855 3135
rect 31855 1159 31864 3135
rect 31908 1159 31917 3135
rect 31917 1159 31951 3135
rect 31951 1159 31960 3135
rect 32004 1159 32013 3135
rect 32013 1159 32047 3135
rect 32047 1159 32056 3135
rect 32100 1159 32109 3135
rect 32109 1159 32143 3135
rect 32143 1159 32152 3135
rect 32196 1159 32205 3135
rect 32205 1159 32239 3135
rect 32239 1159 32248 3135
rect 32292 1159 32301 3135
rect 32301 1159 32335 3135
rect 32335 1159 32344 3135
rect 32388 1159 32397 3135
rect 32397 1159 32431 3135
rect 32431 1159 32440 3135
rect 32484 1159 32493 3135
rect 32493 1159 32527 3135
rect 32527 1159 32536 3135
rect 32580 1159 32589 3135
rect 32589 1159 32623 3135
rect 32623 1159 32632 3135
rect 32676 1159 32685 3135
rect 32685 1159 32719 3135
rect 32719 1159 32728 3135
rect 32772 1159 32781 3135
rect 32781 1159 32815 3135
rect 32815 1159 32824 3135
rect 32868 1159 32877 3135
rect 32877 1159 32911 3135
rect 32911 1159 32920 3135
rect 32964 1159 32973 3135
rect 32973 1159 33007 3135
rect 33007 1159 33016 3135
rect 33060 1159 33069 3135
rect 33069 1159 33103 3135
rect 33103 1159 33112 3135
rect 33156 1159 33165 3135
rect 33165 1159 33199 3135
rect 33199 1159 33208 3135
rect 33252 1159 33261 3135
rect 33261 1159 33295 3135
rect 33295 1159 33304 3135
rect 33348 1159 33357 3135
rect 33357 1159 33391 3135
rect 33391 1159 33400 3135
rect 33444 1159 33453 3135
rect 33453 1159 33487 3135
rect 33487 1159 33496 3135
rect 33540 1159 33549 3135
rect 33549 1159 33583 3135
rect 33583 1159 33592 3135
rect 33636 1159 33645 3135
rect 33645 1159 33679 3135
rect 33679 1159 33688 3135
rect 33732 1159 33741 3135
rect 33741 1159 33775 3135
rect 33775 1159 33784 3135
rect 33828 1159 33837 3135
rect 33837 1159 33871 3135
rect 33871 1159 33880 3135
rect 33924 1159 33933 3135
rect 33933 1159 33967 3135
rect 33967 1159 33976 3135
rect 34020 1159 34029 3135
rect 34029 1159 34063 3135
rect 34063 1159 34072 3135
rect 34116 1159 34125 3135
rect 34125 1159 34159 3135
rect 34159 1159 34168 3135
rect 34212 1159 34221 3135
rect 34221 1159 34255 3135
rect 34255 1159 34264 3135
rect 34308 1159 34317 3135
rect 34317 1159 34351 3135
rect 34351 1159 34360 3135
rect 34404 1159 34413 3135
rect 34413 1159 34447 3135
rect 34447 1159 34456 3135
rect 34500 1159 34509 3135
rect 34509 1159 34543 3135
rect 34543 1159 34552 3135
rect 34596 1159 34605 3135
rect 34605 1159 34639 3135
rect 34639 1159 34648 3135
rect 34692 1159 34701 3135
rect 34701 1159 34735 3135
rect 34735 1159 34744 3135
rect 34788 1159 34797 3135
rect 34797 1159 34831 3135
rect 34831 1159 34840 3135
rect 34884 1159 34893 3135
rect 34893 1159 34927 3135
rect 34927 1159 34936 3135
rect 34980 1159 34989 3135
rect 34989 1159 35023 3135
rect 35023 1159 35032 3135
rect 35076 1159 35085 3135
rect 35085 1159 35119 3135
rect 35119 1159 35128 3135
rect 35172 1159 35181 3135
rect 35181 1159 35215 3135
rect 35215 1159 35224 3135
rect 35268 1159 35277 3135
rect 35277 1159 35311 3135
rect 35311 1159 35320 3135
rect 35364 1159 35373 3135
rect 35373 1159 35407 3135
rect 35407 1159 35416 3135
rect 35460 1159 35469 3135
rect 35469 1159 35503 3135
rect 35503 1159 35512 3135
rect 35556 1159 35565 3135
rect 35565 1159 35599 3135
rect 35599 1159 35608 3135
rect 35652 1159 35661 3135
rect 35661 1159 35695 3135
rect 35695 1159 35704 3135
rect 35748 1159 35757 3135
rect 35757 1159 35791 3135
rect 35791 1159 35800 3135
rect 35844 1159 35853 3135
rect 35853 1159 35887 3135
rect 35887 1159 35896 3135
rect 35940 1159 35949 3135
rect 35949 1159 35983 3135
rect 35983 1159 35992 3135
rect 36036 1159 36045 3135
rect 36045 1159 36079 3135
rect 36079 1159 36088 3135
rect 36132 1159 36141 3135
rect 36141 1159 36175 3135
rect 36175 1159 36184 3135
rect 36228 1159 36237 3135
rect 36237 1159 36271 3135
rect 36271 1159 36280 3135
rect 36324 1159 36333 3135
rect 36333 1159 36367 3135
rect 36367 1159 36376 3135
rect 36420 1159 36429 3135
rect 36429 1159 36463 3135
rect 36463 1159 36472 3135
rect 36516 1159 36525 3135
rect 36525 1159 36559 3135
rect 36559 1159 36568 3135
rect 36612 1159 36621 3135
rect 36621 1159 36655 3135
rect 36655 1159 36664 3135
rect 36708 1159 36717 3135
rect 36717 1159 36751 3135
rect 36751 1159 36760 3135
rect 36804 1159 36813 3135
rect 36813 1159 36847 3135
rect 36847 1159 36856 3135
rect 36900 1159 36909 3135
rect 36909 1159 36943 3135
rect 36943 1159 36952 3135
rect 36996 1159 37005 3135
rect 37005 1159 37039 3135
rect 37039 1159 37048 3135
rect 37092 1159 37101 3135
rect 37101 1159 37135 3135
rect 37135 1159 37144 3135
rect 37188 1159 37197 3135
rect 37197 1159 37231 3135
rect 37231 1159 37240 3135
rect 37284 1159 37293 3135
rect 37293 1159 37327 3135
rect 37327 1159 37336 3135
rect 37380 1159 37389 3135
rect 37389 1159 37423 3135
rect 37423 1159 37432 3135
rect 37476 1159 37485 3135
rect 37485 1159 37519 3135
rect 37519 1159 37528 3135
rect 37572 1159 37581 3135
rect 37581 1159 37615 3135
rect 37615 1159 37624 3135
rect 37668 1159 37677 3135
rect 37677 1159 37711 3135
rect 37711 1159 37720 3135
rect 37764 1159 37773 3135
rect 37773 1159 37807 3135
rect 37807 1159 37816 3135
rect 37860 1159 37869 3135
rect 37869 1159 37903 3135
rect 37903 1159 37912 3135
rect 37956 1159 37965 3135
rect 37965 1159 37999 3135
rect 37999 1159 38008 3135
rect 38052 1159 38061 3135
rect 38061 1159 38095 3135
rect 38095 1159 38104 3135
rect 38148 1159 38157 3135
rect 38157 1159 38191 3135
rect 38191 1159 38200 3135
rect 38244 1159 38253 3135
rect 38253 1159 38287 3135
rect 38287 1159 38296 3135
rect 38340 1159 38349 3135
rect 38349 1159 38383 3135
rect 38383 1159 38392 3135
rect 38436 1159 38445 3135
rect 38445 1159 38479 3135
rect 38479 1159 38488 3135
rect 38532 1159 38541 3135
rect 38541 1159 38575 3135
rect 38575 1159 38584 3135
rect 38628 1158 38637 3134
rect 38637 1158 38671 3134
rect 38671 1158 38680 3134
<< metal2 >>
rect 29025 3135 29083 3147
rect 29025 1159 29028 3135
rect 29080 1159 29083 3135
rect 29025 830 29083 1159
rect 29121 3135 29179 3147
rect 29121 1159 29122 3135
rect 29178 1159 29179 3135
rect 29121 1147 29179 1159
rect 29217 3135 29275 3147
rect 29217 1159 29220 3135
rect 29272 1159 29275 3135
rect 29217 830 29275 1159
rect 29313 3135 29371 3147
rect 29313 1159 29314 3135
rect 29370 1159 29371 3135
rect 29313 1147 29371 1159
rect 29409 3135 29467 3147
rect 29409 1159 29412 3135
rect 29464 1159 29467 3135
rect 29409 830 29467 1159
rect 29505 3135 29563 3147
rect 29505 1159 29506 3135
rect 29562 1159 29563 3135
rect 29505 1147 29563 1159
rect 29601 3135 29659 3147
rect 29601 1159 29604 3135
rect 29656 1159 29659 3135
rect 29601 830 29659 1159
rect 29697 3135 29755 3147
rect 29697 1159 29698 3135
rect 29754 1159 29755 3135
rect 29697 1147 29755 1159
rect 29793 3135 29851 3147
rect 29793 1159 29796 3135
rect 29848 1159 29851 3135
rect 29793 830 29851 1159
rect 29889 3135 29947 3147
rect 29889 1159 29890 3135
rect 29946 1159 29947 3135
rect 29889 1147 29947 1159
rect 29985 3135 30043 3147
rect 29985 1159 29988 3135
rect 30040 1159 30043 3135
rect 29985 830 30043 1159
rect 30081 3135 30139 3147
rect 30081 1159 30082 3135
rect 30138 1159 30139 3135
rect 30081 1147 30139 1159
rect 30177 3135 30235 3147
rect 30177 1159 30180 3135
rect 30232 1159 30235 3135
rect 30177 830 30235 1159
rect 30273 3135 30331 3147
rect 30273 1159 30274 3135
rect 30330 1159 30331 3135
rect 30273 1147 30331 1159
rect 30369 3135 30427 3147
rect 30369 1159 30372 3135
rect 30424 1159 30427 3135
rect 30369 830 30427 1159
rect 30465 3135 30523 3147
rect 30465 1159 30466 3135
rect 30522 1159 30523 3135
rect 30465 1147 30523 1159
rect 30561 3135 30619 3147
rect 30561 1159 30564 3135
rect 30616 1159 30619 3135
rect 30561 830 30619 1159
rect 30657 3135 30715 3147
rect 30657 1159 30658 3135
rect 30714 1159 30715 3135
rect 30657 1147 30715 1159
rect 30753 3135 30811 3147
rect 30753 1159 30756 3135
rect 30808 1159 30811 3135
rect 30753 830 30811 1159
rect 30849 3135 30907 3147
rect 30849 1159 30850 3135
rect 30906 1159 30907 3135
rect 30849 1147 30907 1159
rect 30945 3135 31003 3147
rect 30945 1159 30948 3135
rect 31000 1159 31003 3135
rect 30945 830 31003 1159
rect 31041 3135 31099 3147
rect 31041 1159 31042 3135
rect 31098 1159 31099 3135
rect 31041 1147 31099 1159
rect 31137 3135 31195 3147
rect 31137 1159 31140 3135
rect 31192 1159 31195 3135
rect 31137 830 31195 1159
rect 31233 3135 31291 3147
rect 31233 1159 31234 3135
rect 31290 1159 31291 3135
rect 31233 1147 31291 1159
rect 31329 3135 31387 3147
rect 31329 1159 31332 3135
rect 31384 1159 31387 3135
rect 31329 830 31387 1159
rect 31425 3135 31483 3147
rect 31425 1159 31426 3135
rect 31482 1159 31483 3135
rect 31425 1147 31483 1159
rect 31521 3135 31579 3147
rect 31521 1159 31524 3135
rect 31576 1159 31579 3135
rect 31521 830 31579 1159
rect 31617 3135 31675 3147
rect 31617 1159 31618 3135
rect 31674 1159 31675 3135
rect 31617 1147 31675 1159
rect 31713 3135 31771 3147
rect 31713 1159 31716 3135
rect 31768 1159 31771 3135
rect 31713 830 31771 1159
rect 31809 3135 31867 3147
rect 31809 1159 31810 3135
rect 31866 1159 31867 3135
rect 31809 1147 31867 1159
rect 31905 3135 31963 3147
rect 31905 1159 31908 3135
rect 31960 1159 31963 3135
rect 31905 830 31963 1159
rect 32001 3135 32059 3147
rect 32001 1159 32002 3135
rect 32058 1159 32059 3135
rect 32001 1147 32059 1159
rect 32097 3135 32155 3147
rect 32097 1159 32100 3135
rect 32152 1159 32155 3135
rect 32097 830 32155 1159
rect 32193 3135 32251 3147
rect 32193 1159 32194 3135
rect 32250 1159 32251 3135
rect 32193 1147 32251 1159
rect 32289 3135 32347 3147
rect 32289 1159 32292 3135
rect 32344 1159 32347 3135
rect 32289 830 32347 1159
rect 32385 3135 32443 3147
rect 32385 1159 32386 3135
rect 32442 1159 32443 3135
rect 32385 1147 32443 1159
rect 32481 3135 32539 3147
rect 32481 1159 32484 3135
rect 32536 1159 32539 3135
rect 32481 830 32539 1159
rect 32577 3135 32635 3147
rect 32577 1159 32578 3135
rect 32634 1159 32635 3135
rect 32577 1147 32635 1159
rect 32673 3135 32731 3147
rect 32673 1159 32676 3135
rect 32728 1159 32731 3135
rect 32673 830 32731 1159
rect 32769 3135 32827 3147
rect 32769 1159 32770 3135
rect 32826 1159 32827 3135
rect 32769 1147 32827 1159
rect 32865 3135 32923 3147
rect 32865 1159 32868 3135
rect 32920 1159 32923 3135
rect 32865 830 32923 1159
rect 32961 3135 33019 3147
rect 32961 1159 32962 3135
rect 33018 1159 33019 3135
rect 32961 1147 33019 1159
rect 33057 3135 33115 3147
rect 33057 1159 33060 3135
rect 33112 1159 33115 3135
rect 33057 830 33115 1159
rect 33153 3135 33211 3147
rect 33153 1159 33154 3135
rect 33210 1159 33211 3135
rect 33153 1147 33211 1159
rect 33249 3135 33307 3147
rect 33249 1159 33252 3135
rect 33304 1159 33307 3135
rect 33249 830 33307 1159
rect 33345 3135 33403 3147
rect 33345 1159 33346 3135
rect 33402 1159 33403 3135
rect 33345 1147 33403 1159
rect 33441 3135 33499 3147
rect 33441 1159 33444 3135
rect 33496 1159 33499 3135
rect 33441 830 33499 1159
rect 33537 3135 33595 3147
rect 33537 1159 33538 3135
rect 33594 1159 33595 3135
rect 33537 1147 33595 1159
rect 33633 3135 33691 3147
rect 33633 1159 33636 3135
rect 33688 1159 33691 3135
rect 33633 830 33691 1159
rect 33729 3135 33787 3147
rect 33729 1159 33730 3135
rect 33786 1159 33787 3135
rect 33729 1147 33787 1159
rect 33825 3135 33883 3147
rect 33825 1159 33828 3135
rect 33880 1159 33883 3135
rect 33825 830 33883 1159
rect 33921 3135 33979 3147
rect 33921 1159 33922 3135
rect 33978 1159 33979 3135
rect 33921 1147 33979 1159
rect 34017 3135 34075 3147
rect 34017 1159 34020 3135
rect 34072 1159 34075 3135
rect 34017 830 34075 1159
rect 34113 3135 34171 3147
rect 34113 1159 34114 3135
rect 34170 1159 34171 3135
rect 34113 1147 34171 1159
rect 34209 3135 34267 3147
rect 34209 1159 34212 3135
rect 34264 1159 34267 3135
rect 34209 830 34267 1159
rect 34305 3135 34363 3147
rect 34305 1159 34306 3135
rect 34362 1159 34363 3135
rect 34305 1147 34363 1159
rect 34401 3135 34459 3147
rect 34401 1159 34404 3135
rect 34456 1159 34459 3135
rect 34401 830 34459 1159
rect 34497 3135 34555 3147
rect 34497 1159 34498 3135
rect 34554 1159 34555 3135
rect 34497 1147 34555 1159
rect 34593 3135 34651 3147
rect 34593 1159 34596 3135
rect 34648 1159 34651 3135
rect 34593 830 34651 1159
rect 34689 3135 34747 3147
rect 34689 1159 34690 3135
rect 34746 1159 34747 3135
rect 34689 1147 34747 1159
rect 34785 3135 34843 3147
rect 34785 1159 34788 3135
rect 34840 1159 34843 3135
rect 34785 830 34843 1159
rect 34881 3135 34939 3147
rect 34881 1159 34882 3135
rect 34938 1159 34939 3135
rect 34881 1147 34939 1159
rect 34977 3135 35035 3147
rect 34977 1159 34980 3135
rect 35032 1159 35035 3135
rect 34977 830 35035 1159
rect 35073 3135 35131 3147
rect 35073 1159 35074 3135
rect 35130 1159 35131 3135
rect 35073 1147 35131 1159
rect 35169 3135 35227 3147
rect 35169 1159 35172 3135
rect 35224 1159 35227 3135
rect 35169 830 35227 1159
rect 35265 3135 35323 3147
rect 35265 1159 35266 3135
rect 35322 1159 35323 3135
rect 35265 1147 35323 1159
rect 35361 3135 35419 3147
rect 35361 1159 35364 3135
rect 35416 1159 35419 3135
rect 35361 830 35419 1159
rect 35457 3135 35515 3147
rect 35457 1159 35458 3135
rect 35514 1159 35515 3135
rect 35457 1147 35515 1159
rect 35553 3135 35611 3147
rect 35553 1159 35556 3135
rect 35608 1159 35611 3135
rect 35553 830 35611 1159
rect 35649 3135 35707 3147
rect 35649 1159 35650 3135
rect 35706 1159 35707 3135
rect 35649 1147 35707 1159
rect 35745 3135 35803 3147
rect 35745 1159 35748 3135
rect 35800 1159 35803 3135
rect 35745 830 35803 1159
rect 35841 3135 35899 3147
rect 35841 1159 35842 3135
rect 35898 1159 35899 3135
rect 35841 1147 35899 1159
rect 35937 3135 35995 3147
rect 35937 1159 35940 3135
rect 35992 1159 35995 3135
rect 35937 830 35995 1159
rect 36033 3135 36091 3147
rect 36033 1159 36034 3135
rect 36090 1159 36091 3135
rect 36033 1147 36091 1159
rect 36129 3135 36187 3147
rect 36129 1159 36132 3135
rect 36184 1159 36187 3135
rect 36129 830 36187 1159
rect 36225 3135 36283 3147
rect 36225 1159 36226 3135
rect 36282 1159 36283 3135
rect 36225 1147 36283 1159
rect 36321 3135 36379 3147
rect 36321 1159 36324 3135
rect 36376 1159 36379 3135
rect 36321 830 36379 1159
rect 36417 3135 36475 3147
rect 36417 1159 36418 3135
rect 36474 1159 36475 3135
rect 36417 1147 36475 1159
rect 36513 3135 36571 3147
rect 36513 1159 36516 3135
rect 36568 1159 36571 3135
rect 36513 830 36571 1159
rect 36609 3135 36667 3147
rect 36609 1159 36610 3135
rect 36666 1159 36667 3135
rect 36609 1147 36667 1159
rect 36705 3135 36763 3147
rect 36705 1159 36708 3135
rect 36760 1159 36763 3135
rect 36705 830 36763 1159
rect 36801 3135 36859 3147
rect 36801 1159 36802 3135
rect 36858 1159 36859 3135
rect 36801 1147 36859 1159
rect 36897 3135 36955 3147
rect 36897 1159 36900 3135
rect 36952 1159 36955 3135
rect 36897 830 36955 1159
rect 36993 3135 37051 3147
rect 36993 1159 36994 3135
rect 37050 1159 37051 3135
rect 36993 1147 37051 1159
rect 37089 3135 37147 3147
rect 37089 1159 37092 3135
rect 37144 1159 37147 3135
rect 37089 830 37147 1159
rect 37185 3135 37243 3147
rect 37185 1159 37186 3135
rect 37242 1159 37243 3135
rect 37185 1147 37243 1159
rect 37281 3135 37339 3147
rect 37281 1159 37284 3135
rect 37336 1159 37339 3135
rect 37281 830 37339 1159
rect 37377 3135 37435 3147
rect 37377 1159 37378 3135
rect 37434 1159 37435 3135
rect 37377 1147 37435 1159
rect 37473 3135 37531 3147
rect 37473 1159 37476 3135
rect 37528 1159 37531 3135
rect 37473 830 37531 1159
rect 37569 3135 37627 3147
rect 37569 1159 37570 3135
rect 37626 1159 37627 3135
rect 37569 1147 37627 1159
rect 37665 3135 37723 3147
rect 37665 1159 37668 3135
rect 37720 1159 37723 3135
rect 37665 830 37723 1159
rect 37761 3135 37819 3147
rect 37761 1159 37762 3135
rect 37818 1159 37819 3135
rect 37761 1147 37819 1159
rect 37857 3135 37915 3147
rect 37857 1159 37860 3135
rect 37912 1159 37915 3135
rect 37857 830 37915 1159
rect 37953 3135 38011 3147
rect 37953 1159 37954 3135
rect 38010 1159 38011 3135
rect 37953 1147 38011 1159
rect 38049 3135 38107 3147
rect 38049 1159 38052 3135
rect 38104 1159 38107 3135
rect 38049 830 38107 1159
rect 38145 3135 38203 3147
rect 38145 1159 38146 3135
rect 38202 1159 38203 3135
rect 38145 1147 38203 1159
rect 38241 3135 38299 3147
rect 38241 1159 38244 3135
rect 38296 1159 38299 3135
rect 38241 830 38299 1159
rect 38337 3135 38395 3147
rect 38337 1159 38338 3135
rect 38394 1159 38395 3135
rect 38337 1147 38395 1159
rect 38433 3135 38491 3147
rect 38433 1159 38436 3135
rect 38488 1159 38491 3135
rect 38433 830 38491 1159
rect 38529 3135 38587 3147
rect 38529 1159 38530 3135
rect 38586 1159 38587 3135
rect 38529 1147 38587 1159
rect 38625 3134 38683 3146
rect 38625 1158 38628 3134
rect 38680 1158 38683 3134
rect 38625 830 38683 1158
rect 29025 746 38684 830
rect 38625 745 38683 746
<< via2 >>
rect 29122 1159 29124 3135
rect 29124 1159 29176 3135
rect 29176 1159 29178 3135
rect 29314 1159 29316 3135
rect 29316 1159 29368 3135
rect 29368 1159 29370 3135
rect 29506 1159 29508 3135
rect 29508 1159 29560 3135
rect 29560 1159 29562 3135
rect 29698 1159 29700 3135
rect 29700 1159 29752 3135
rect 29752 1159 29754 3135
rect 29890 1159 29892 3135
rect 29892 1159 29944 3135
rect 29944 1159 29946 3135
rect 30082 1159 30084 3135
rect 30084 1159 30136 3135
rect 30136 1159 30138 3135
rect 30274 1159 30276 3135
rect 30276 1159 30328 3135
rect 30328 1159 30330 3135
rect 30466 1159 30468 3135
rect 30468 1159 30520 3135
rect 30520 1159 30522 3135
rect 30658 1159 30660 3135
rect 30660 1159 30712 3135
rect 30712 1159 30714 3135
rect 30850 1159 30852 3135
rect 30852 1159 30904 3135
rect 30904 1159 30906 3135
rect 31042 1159 31044 3135
rect 31044 1159 31096 3135
rect 31096 1159 31098 3135
rect 31234 1159 31236 3135
rect 31236 1159 31288 3135
rect 31288 1159 31290 3135
rect 31426 1159 31428 3135
rect 31428 1159 31480 3135
rect 31480 1159 31482 3135
rect 31618 1159 31620 3135
rect 31620 1159 31672 3135
rect 31672 1159 31674 3135
rect 31810 1159 31812 3135
rect 31812 1159 31864 3135
rect 31864 1159 31866 3135
rect 32002 1159 32004 3135
rect 32004 1159 32056 3135
rect 32056 1159 32058 3135
rect 32194 1159 32196 3135
rect 32196 1159 32248 3135
rect 32248 1159 32250 3135
rect 32386 1159 32388 3135
rect 32388 1159 32440 3135
rect 32440 1159 32442 3135
rect 32578 1159 32580 3135
rect 32580 1159 32632 3135
rect 32632 1159 32634 3135
rect 32770 1159 32772 3135
rect 32772 1159 32824 3135
rect 32824 1159 32826 3135
rect 32962 1159 32964 3135
rect 32964 1159 33016 3135
rect 33016 1159 33018 3135
rect 33154 1159 33156 3135
rect 33156 1159 33208 3135
rect 33208 1159 33210 3135
rect 33346 1159 33348 3135
rect 33348 1159 33400 3135
rect 33400 1159 33402 3135
rect 33538 1159 33540 3135
rect 33540 1159 33592 3135
rect 33592 1159 33594 3135
rect 33730 1159 33732 3135
rect 33732 1159 33784 3135
rect 33784 1159 33786 3135
rect 33922 1159 33924 3135
rect 33924 1159 33976 3135
rect 33976 1159 33978 3135
rect 34114 1159 34116 3135
rect 34116 1159 34168 3135
rect 34168 1159 34170 3135
rect 34306 1159 34308 3135
rect 34308 1159 34360 3135
rect 34360 1159 34362 3135
rect 34498 1159 34500 3135
rect 34500 1159 34552 3135
rect 34552 1159 34554 3135
rect 34690 1159 34692 3135
rect 34692 1159 34744 3135
rect 34744 1159 34746 3135
rect 34882 1159 34884 3135
rect 34884 1159 34936 3135
rect 34936 1159 34938 3135
rect 35074 1159 35076 3135
rect 35076 1159 35128 3135
rect 35128 1159 35130 3135
rect 35266 1159 35268 3135
rect 35268 1159 35320 3135
rect 35320 1159 35322 3135
rect 35458 1159 35460 3135
rect 35460 1159 35512 3135
rect 35512 1159 35514 3135
rect 35650 1159 35652 3135
rect 35652 1159 35704 3135
rect 35704 1159 35706 3135
rect 35842 1159 35844 3135
rect 35844 1159 35896 3135
rect 35896 1159 35898 3135
rect 36034 1159 36036 3135
rect 36036 1159 36088 3135
rect 36088 1159 36090 3135
rect 36226 1159 36228 3135
rect 36228 1159 36280 3135
rect 36280 1159 36282 3135
rect 36418 1159 36420 3135
rect 36420 1159 36472 3135
rect 36472 1159 36474 3135
rect 36610 1159 36612 3135
rect 36612 1159 36664 3135
rect 36664 1159 36666 3135
rect 36802 1159 36804 3135
rect 36804 1159 36856 3135
rect 36856 1159 36858 3135
rect 36994 1159 36996 3135
rect 36996 1159 37048 3135
rect 37048 1159 37050 3135
rect 37186 1159 37188 3135
rect 37188 1159 37240 3135
rect 37240 1159 37242 3135
rect 37378 1159 37380 3135
rect 37380 1159 37432 3135
rect 37432 1159 37434 3135
rect 37570 1159 37572 3135
rect 37572 1159 37624 3135
rect 37624 1159 37626 3135
rect 37762 1159 37764 3135
rect 37764 1159 37816 3135
rect 37816 1159 37818 3135
rect 37954 1159 37956 3135
rect 37956 1159 38008 3135
rect 38008 1159 38010 3135
rect 38146 1159 38148 3135
rect 38148 1159 38200 3135
rect 38200 1159 38202 3135
rect 38338 1159 38340 3135
rect 38340 1159 38392 3135
rect 38392 1159 38394 3135
rect 38530 1159 38532 3135
rect 38532 1159 38584 3135
rect 38584 1159 38586 3135
<< metal3 >>
rect 29116 3522 38592 3606
rect 29116 3135 29184 3522
rect 29116 1159 29122 3135
rect 29178 1159 29184 3135
rect 29116 1147 29184 1159
rect 29308 3135 29376 3522
rect 29308 1159 29314 3135
rect 29370 1159 29376 3135
rect 29308 1147 29376 1159
rect 29500 3135 29568 3522
rect 29500 1159 29506 3135
rect 29562 1159 29568 3135
rect 29500 1147 29568 1159
rect 29692 3135 29760 3522
rect 29692 1159 29698 3135
rect 29754 1159 29760 3135
rect 29692 1147 29760 1159
rect 29884 3135 29952 3522
rect 29884 1159 29890 3135
rect 29946 1159 29952 3135
rect 29884 1147 29952 1159
rect 30076 3135 30144 3522
rect 30076 1159 30082 3135
rect 30138 1159 30144 3135
rect 30076 1147 30144 1159
rect 30268 3135 30336 3522
rect 30268 1159 30274 3135
rect 30330 1159 30336 3135
rect 30268 1147 30336 1159
rect 30460 3135 30528 3522
rect 30460 1159 30466 3135
rect 30522 1159 30528 3135
rect 30460 1147 30528 1159
rect 30652 3135 30720 3522
rect 30652 1159 30658 3135
rect 30714 1159 30720 3135
rect 30652 1147 30720 1159
rect 30844 3135 30912 3522
rect 30844 1159 30850 3135
rect 30906 1159 30912 3135
rect 30844 1147 30912 1159
rect 31036 3135 31104 3522
rect 31036 1159 31042 3135
rect 31098 1159 31104 3135
rect 31036 1147 31104 1159
rect 31228 3135 31296 3522
rect 31228 1159 31234 3135
rect 31290 1159 31296 3135
rect 31228 1147 31296 1159
rect 31420 3135 31488 3522
rect 31420 1159 31426 3135
rect 31482 1159 31488 3135
rect 31420 1147 31488 1159
rect 31612 3135 31680 3522
rect 31612 1159 31618 3135
rect 31674 1159 31680 3135
rect 31612 1147 31680 1159
rect 31804 3135 31872 3522
rect 31804 1159 31810 3135
rect 31866 1159 31872 3135
rect 31804 1147 31872 1159
rect 31996 3135 32064 3522
rect 31996 1159 32002 3135
rect 32058 1159 32064 3135
rect 31996 1147 32064 1159
rect 32188 3135 32256 3522
rect 32188 1159 32194 3135
rect 32250 1159 32256 3135
rect 32188 1147 32256 1159
rect 32380 3135 32448 3522
rect 32380 1159 32386 3135
rect 32442 1159 32448 3135
rect 32380 1147 32448 1159
rect 32572 3135 32640 3522
rect 32572 1159 32578 3135
rect 32634 1159 32640 3135
rect 32572 1147 32640 1159
rect 32764 3135 32832 3522
rect 32764 1159 32770 3135
rect 32826 1159 32832 3135
rect 32764 1147 32832 1159
rect 32956 3135 33024 3522
rect 32956 1159 32962 3135
rect 33018 1159 33024 3135
rect 32956 1147 33024 1159
rect 33148 3135 33216 3522
rect 33148 1159 33154 3135
rect 33210 1159 33216 3135
rect 33148 1147 33216 1159
rect 33340 3135 33408 3522
rect 33340 1159 33346 3135
rect 33402 1159 33408 3135
rect 33340 1147 33408 1159
rect 33532 3135 33600 3522
rect 33532 1159 33538 3135
rect 33594 1159 33600 3135
rect 33532 1147 33600 1159
rect 33724 3135 33792 3522
rect 33724 1159 33730 3135
rect 33786 1159 33792 3135
rect 33724 1147 33792 1159
rect 33916 3135 33984 3522
rect 33916 1159 33922 3135
rect 33978 1159 33984 3135
rect 33916 1147 33984 1159
rect 34108 3135 34176 3522
rect 34108 1159 34114 3135
rect 34170 1159 34176 3135
rect 34108 1147 34176 1159
rect 34300 3135 34368 3522
rect 34300 1159 34306 3135
rect 34362 1159 34368 3135
rect 34300 1147 34368 1159
rect 34492 3135 34560 3522
rect 34492 1159 34498 3135
rect 34554 1159 34560 3135
rect 34492 1147 34560 1159
rect 34684 3135 34752 3522
rect 34684 1159 34690 3135
rect 34746 1159 34752 3135
rect 34684 1147 34752 1159
rect 34876 3135 34944 3522
rect 34876 1159 34882 3135
rect 34938 1159 34944 3135
rect 34876 1147 34944 1159
rect 35068 3135 35136 3522
rect 35068 1159 35074 3135
rect 35130 1159 35136 3135
rect 35068 1147 35136 1159
rect 35260 3135 35328 3522
rect 35260 1159 35266 3135
rect 35322 1159 35328 3135
rect 35260 1147 35328 1159
rect 35452 3135 35520 3522
rect 35452 1159 35458 3135
rect 35514 1159 35520 3135
rect 35452 1147 35520 1159
rect 35644 3135 35712 3522
rect 35644 1159 35650 3135
rect 35706 1159 35712 3135
rect 35644 1147 35712 1159
rect 35836 3135 35904 3522
rect 35836 1159 35842 3135
rect 35898 1159 35904 3135
rect 35836 1147 35904 1159
rect 36028 3135 36096 3522
rect 36028 1159 36034 3135
rect 36090 1159 36096 3135
rect 36028 1147 36096 1159
rect 36220 3135 36288 3522
rect 36220 1159 36226 3135
rect 36282 1159 36288 3135
rect 36220 1147 36288 1159
rect 36412 3135 36480 3522
rect 36412 1159 36418 3135
rect 36474 1159 36480 3135
rect 36412 1147 36480 1159
rect 36604 3135 36672 3522
rect 36604 1159 36610 3135
rect 36666 1159 36672 3135
rect 36604 1147 36672 1159
rect 36796 3135 36864 3522
rect 36796 1159 36802 3135
rect 36858 1159 36864 3135
rect 36796 1147 36864 1159
rect 36988 3135 37056 3522
rect 36988 1159 36994 3135
rect 37050 1159 37056 3135
rect 36988 1147 37056 1159
rect 37180 3135 37248 3522
rect 37180 1159 37186 3135
rect 37242 1159 37248 3135
rect 37180 1147 37248 1159
rect 37372 3135 37440 3522
rect 37372 1159 37378 3135
rect 37434 1159 37440 3135
rect 37372 1147 37440 1159
rect 37564 3135 37632 3522
rect 37564 1159 37570 3135
rect 37626 1159 37632 3135
rect 37564 1147 37632 1159
rect 37756 3135 37824 3522
rect 37756 1159 37762 3135
rect 37818 1159 37824 3135
rect 37756 1147 37824 1159
rect 37948 3135 38016 3522
rect 37948 1159 37954 3135
rect 38010 1159 38016 3135
rect 37948 1147 38016 1159
rect 38140 3135 38208 3522
rect 38140 1159 38146 3135
rect 38202 1159 38208 3135
rect 38140 1147 38208 1159
rect 38332 3135 38400 3522
rect 38332 1159 38338 3135
rect 38394 1159 38400 3135
rect 38332 1147 38400 1159
rect 38524 3135 38592 3522
rect 38524 1159 38530 3135
rect 38586 1159 38592 3135
rect 38524 1147 38592 1159
use sky130_fd_pr__nfet_01v8_spf0jm  sky130_fd_pr__nfet_01v8_spf0jm_0
timestamp 1606421359
transform 1 0 33854 0 1 2147
box -4967 -1210 4967 1210
<< end >>
